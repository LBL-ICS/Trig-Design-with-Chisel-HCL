module VCORDIC(
  input         clock,
  input         reset,
  input  [31:0] io_in_y0,
  output [31:0] io_out_z
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] tofixedx0_io_in; // @[VCORDIC.scala 107:33]
  wire [63:0] tofixedx0_io_out; // @[VCORDIC.scala 107:33]
  wire [31:0] tofixedy0_io_in; // @[VCORDIC.scala 108:33]
  wire [63:0] tofixedy0_io_out; // @[VCORDIC.scala 108:33]
  wire [31:0] tofixedz0_io_in; // @[VCORDIC.scala 109:33]
  wire [63:0] tofixedz0_io_out; // @[VCORDIC.scala 109:33]
  wire [63:0] tofloatxout_io_in; // @[VCORDIC.scala 467:29]
  wire [31:0] tofloatxout_io_out; // @[VCORDIC.scala 467:29]
  wire [63:0] tofloatyout_io_in; // @[VCORDIC.scala 468:29]
  wire [31:0] tofloatyout_io_out; // @[VCORDIC.scala 468:29]
  wire [63:0] tofloatzout_io_in; // @[VCORDIC.scala 469:29]
  wire [31:0] tofloatzout_io_out; // @[VCORDIC.scala 469:29]
  reg [63:0] xr_0; // @[VCORDIC.scala 120:27]
  reg [63:0] xr_1; // @[VCORDIC.scala 120:27]
  reg [63:0] yr_0; // @[VCORDIC.scala 121:27]
  reg [63:0] yr_1; // @[VCORDIC.scala 121:27]
  reg [63:0] zr_0; // @[VCORDIC.scala 122:27]
  reg [63:0] zr_1; // @[VCORDIC.scala 122:27]
  wire  _fxxterm_T = $signed(yr_0) < 64'sh0; // @[VCORDIC.scala 424:33]
  wire [63:0] _fxxterm_T_3 = 64'sh0 - $signed(xr_0); // @[VCORDIC.scala 424:46]
  wire [63:0] fxxterm = $signed(yr_0) < 64'sh0 ? $signed(_fxxterm_T_3) : $signed(xr_0); // @[VCORDIC.scala 424:26]
  wire [63:0] _fxyterm_T_3 = 64'sh0 - $signed(yr_0); // @[VCORDIC.scala 425:46]
  wire [63:0] fxyterm = _fxxterm_T ? $signed(_fxyterm_T_3) : $signed(yr_0); // @[VCORDIC.scala 425:26]
  wire [63:0] _fxthetaterm_T_2 = 64'h0 - 64'hc90fdb00; // @[VCORDIC.scala 426:50]
  wire [63:0] x_1 = $signed(xr_0) + $signed(fxyterm); // @[VCORDIC.scala 428:27]
  wire [63:0] y_1 = $signed(yr_0) - $signed(fxxterm); // @[VCORDIC.scala 429:27]
  wire [63:0] _z_1_T = _fxxterm_T ? _fxthetaterm_T_2 : 64'hc90fdb00; // @[VCORDIC.scala 430:41]
  wire [63:0] z_1 = $signed(zr_0) + $signed(_z_1_T); // @[VCORDIC.scala 430:27]
  wire  _fxxterm_T_4 = $signed(y_1) < 64'sh0; // @[VCORDIC.scala 454:32]
  wire [63:0] _fxxterm_T_7 = 64'sh0 - $signed(x_1); // @[VCORDIC.scala 454:45]
  wire [63:0] fxxterm_1 = $signed(y_1) < 64'sh0 ? $signed(_fxxterm_T_7) : $signed(x_1); // @[VCORDIC.scala 454:26]
  wire [63:0] _fxyterm_T_7 = 64'sh0 - $signed(y_1); // @[VCORDIC.scala 455:45]
  wire [63:0] fxyterm_1 = _fxxterm_T_4 ? $signed(_fxyterm_T_7) : $signed(y_1); // @[VCORDIC.scala 455:26]
  wire [63:0] _fxthetaterm_T_5 = 64'h0 - 64'h76b19c00; // @[VCORDIC.scala 456:49]
  wire [62:0] _GEN_0 = fxyterm_1[63:1]; // @[VCORDIC.scala 458:37]
  wire [63:0] _x_2_T = {{1{_GEN_0[62]}},_GEN_0}; // @[VCORDIC.scala 458:37]
  wire [63:0] x_2 = $signed(x_1) + $signed(_x_2_T); // @[VCORDIC.scala 458:26]
  wire [62:0] _GEN_1 = fxxterm_1[63:1]; // @[VCORDIC.scala 459:37]
  wire [63:0] _y_2_T = {{1{_GEN_1[62]}},_GEN_1}; // @[VCORDIC.scala 459:37]
  wire [63:0] y_2 = $signed(y_1) - $signed(_y_2_T); // @[VCORDIC.scala 459:26]
  wire [63:0] _z_2_T = _fxxterm_T_4 ? _fxthetaterm_T_5 : 64'h76b19c00; // @[VCORDIC.scala 460:40]
  wire [63:0] z_2 = $signed(z_1) + $signed(_z_2_T); // @[VCORDIC.scala 460:26]
  wire  _fxxterm_T_8 = $signed(y_2) < 64'sh0; // @[VCORDIC.scala 454:32]
  wire [63:0] _fxxterm_T_11 = 64'sh0 - $signed(x_2); // @[VCORDIC.scala 454:45]
  wire [63:0] fxxterm_2 = $signed(y_2) < 64'sh0 ? $signed(_fxxterm_T_11) : $signed(x_2); // @[VCORDIC.scala 454:26]
  wire [63:0] _fxyterm_T_11 = 64'sh0 - $signed(y_2); // @[VCORDIC.scala 455:45]
  wire [63:0] fxyterm_2 = _fxxterm_T_8 ? $signed(_fxyterm_T_11) : $signed(y_2); // @[VCORDIC.scala 455:26]
  wire [63:0] _fxthetaterm_T_8 = 64'h0 - 64'h3eb6ec00; // @[VCORDIC.scala 456:49]
  wire [61:0] _GEN_2 = fxyterm_2[63:2]; // @[VCORDIC.scala 458:37]
  wire [63:0] _x_3_T = {{2{_GEN_2[61]}},_GEN_2}; // @[VCORDIC.scala 458:37]
  wire [63:0] x_3 = $signed(x_2) + $signed(_x_3_T); // @[VCORDIC.scala 458:26]
  wire [61:0] _GEN_3 = fxxterm_2[63:2]; // @[VCORDIC.scala 459:37]
  wire [63:0] _y_3_T = {{2{_GEN_3[61]}},_GEN_3}; // @[VCORDIC.scala 459:37]
  wire [63:0] y_3 = $signed(y_2) - $signed(_y_3_T); // @[VCORDIC.scala 459:26]
  wire [63:0] _z_3_T = _fxxterm_T_8 ? _fxthetaterm_T_8 : 64'h3eb6ec00; // @[VCORDIC.scala 460:40]
  wire [63:0] z_3 = $signed(z_2) + $signed(_z_3_T); // @[VCORDIC.scala 460:26]
  wire  _fxxterm_T_12 = $signed(y_3) < 64'sh0; // @[VCORDIC.scala 454:32]
  wire [63:0] _fxxterm_T_15 = 64'sh0 - $signed(x_3); // @[VCORDIC.scala 454:45]
  wire [63:0] fxxterm_3 = $signed(y_3) < 64'sh0 ? $signed(_fxxterm_T_15) : $signed(x_3); // @[VCORDIC.scala 454:26]
  wire [63:0] _fxyterm_T_15 = 64'sh0 - $signed(y_3); // @[VCORDIC.scala 455:45]
  wire [63:0] fxyterm_3 = _fxxterm_T_12 ? $signed(_fxyterm_T_15) : $signed(y_3); // @[VCORDIC.scala 455:26]
  wire [63:0] _fxthetaterm_T_11 = 64'h0 - 64'h1fd5baa0; // @[VCORDIC.scala 456:49]
  wire [60:0] _GEN_4 = fxyterm_3[63:3]; // @[VCORDIC.scala 458:37]
  wire [63:0] _x_4_T = {{3{_GEN_4[60]}},_GEN_4}; // @[VCORDIC.scala 458:37]
  wire [63:0] x_4 = $signed(x_3) + $signed(_x_4_T); // @[VCORDIC.scala 458:26]
  wire [60:0] _GEN_5 = fxxterm_3[63:3]; // @[VCORDIC.scala 459:37]
  wire [63:0] _y_4_T = {{3{_GEN_5[60]}},_GEN_5}; // @[VCORDIC.scala 459:37]
  wire [63:0] y_4 = $signed(y_3) - $signed(_y_4_T); // @[VCORDIC.scala 459:26]
  wire [63:0] _z_4_T = _fxxterm_T_12 ? _fxthetaterm_T_11 : 64'h1fd5baa0; // @[VCORDIC.scala 460:40]
  wire [63:0] z_4 = $signed(z_3) + $signed(_z_4_T); // @[VCORDIC.scala 460:26]
  wire  _fxxterm_T_16 = $signed(y_4) < 64'sh0; // @[VCORDIC.scala 454:32]
  wire [63:0] _fxxterm_T_19 = 64'sh0 - $signed(x_4); // @[VCORDIC.scala 454:45]
  wire [63:0] fxxterm_4 = $signed(y_4) < 64'sh0 ? $signed(_fxxterm_T_19) : $signed(x_4); // @[VCORDIC.scala 454:26]
  wire [63:0] _fxyterm_T_19 = 64'sh0 - $signed(y_4); // @[VCORDIC.scala 455:45]
  wire [63:0] fxyterm_4 = _fxxterm_T_16 ? $signed(_fxyterm_T_19) : $signed(y_4); // @[VCORDIC.scala 455:26]
  wire [63:0] _fxthetaterm_T_14 = 64'h0 - 64'hffaade0; // @[VCORDIC.scala 456:49]
  wire [59:0] _GEN_6 = fxyterm_4[63:4]; // @[VCORDIC.scala 458:37]
  wire [63:0] _x_5_T = {{4{_GEN_6[59]}},_GEN_6}; // @[VCORDIC.scala 458:37]
  wire [63:0] x_5 = $signed(x_4) + $signed(_x_5_T); // @[VCORDIC.scala 458:26]
  wire [59:0] _GEN_7 = fxxterm_4[63:4]; // @[VCORDIC.scala 459:37]
  wire [63:0] _y_5_T = {{4{_GEN_7[59]}},_GEN_7}; // @[VCORDIC.scala 459:37]
  wire [63:0] y_5 = $signed(y_4) - $signed(_y_5_T); // @[VCORDIC.scala 459:26]
  wire [63:0] _z_5_T = _fxxterm_T_16 ? _fxthetaterm_T_14 : 64'hffaade0; // @[VCORDIC.scala 460:40]
  wire [63:0] z_5 = $signed(z_4) + $signed(_z_5_T); // @[VCORDIC.scala 460:26]
  wire  _fxxterm_T_20 = $signed(y_5) < 64'sh0; // @[VCORDIC.scala 454:32]
  wire [63:0] _fxxterm_T_23 = 64'sh0 - $signed(x_5); // @[VCORDIC.scala 454:45]
  wire [63:0] fxxterm_5 = $signed(y_5) < 64'sh0 ? $signed(_fxxterm_T_23) : $signed(x_5); // @[VCORDIC.scala 454:26]
  wire [63:0] _fxyterm_T_23 = 64'sh0 - $signed(y_5); // @[VCORDIC.scala 455:45]
  wire [63:0] fxyterm_5 = _fxxterm_T_20 ? $signed(_fxyterm_T_23) : $signed(y_5); // @[VCORDIC.scala 455:26]
  wire [63:0] _fxthetaterm_T_17 = 64'h0 - 64'h7ff5570; // @[VCORDIC.scala 456:49]
  wire [58:0] _GEN_8 = fxyterm_5[63:5]; // @[VCORDIC.scala 458:37]
  wire [63:0] _x_6_T = {{5{_GEN_8[58]}},_GEN_8}; // @[VCORDIC.scala 458:37]
  wire [63:0] x_6 = $signed(x_5) + $signed(_x_6_T); // @[VCORDIC.scala 458:26]
  wire [58:0] _GEN_9 = fxxterm_5[63:5]; // @[VCORDIC.scala 459:37]
  wire [63:0] _y_6_T = {{5{_GEN_9[58]}},_GEN_9}; // @[VCORDIC.scala 459:37]
  wire [63:0] y_6 = $signed(y_5) - $signed(_y_6_T); // @[VCORDIC.scala 459:26]
  wire [63:0] _z_6_T = _fxxterm_T_20 ? _fxthetaterm_T_17 : 64'h7ff5570; // @[VCORDIC.scala 460:40]
  wire [63:0] z_6 = $signed(z_5) + $signed(_z_6_T); // @[VCORDIC.scala 460:26]
  wire  _fxxterm_T_24 = $signed(y_6) < 64'sh0; // @[VCORDIC.scala 454:32]
  wire [63:0] _fxxterm_T_27 = 64'sh0 - $signed(x_6); // @[VCORDIC.scala 454:45]
  wire [63:0] fxxterm_6 = $signed(y_6) < 64'sh0 ? $signed(_fxxterm_T_27) : $signed(x_6); // @[VCORDIC.scala 454:26]
  wire [63:0] _fxyterm_T_27 = 64'sh0 - $signed(y_6); // @[VCORDIC.scala 455:45]
  wire [63:0] fxyterm_6 = _fxxterm_T_24 ? $signed(_fxyterm_T_27) : $signed(y_6); // @[VCORDIC.scala 455:26]
  wire [63:0] _fxthetaterm_T_20 = 64'h0 - 64'h3ffeaac; // @[VCORDIC.scala 456:49]
  wire [57:0] _GEN_10 = fxyterm_6[63:6]; // @[VCORDIC.scala 458:37]
  wire [63:0] _x_7_T = {{6{_GEN_10[57]}},_GEN_10}; // @[VCORDIC.scala 458:37]
  wire [63:0] x_7 = $signed(x_6) + $signed(_x_7_T); // @[VCORDIC.scala 458:26]
  wire [57:0] _GEN_11 = fxxterm_6[63:6]; // @[VCORDIC.scala 459:37]
  wire [63:0] _y_7_T = {{6{_GEN_11[57]}},_GEN_11}; // @[VCORDIC.scala 459:37]
  wire [63:0] y_7 = $signed(y_6) - $signed(_y_7_T); // @[VCORDIC.scala 459:26]
  wire [63:0] _z_7_T = _fxxterm_T_24 ? _fxthetaterm_T_20 : 64'h3ffeaac; // @[VCORDIC.scala 460:40]
  wire [63:0] z_7 = $signed(z_6) + $signed(_z_7_T); // @[VCORDIC.scala 460:26]
  wire  _fxxterm_T_28 = $signed(y_7) < 64'sh0; // @[VCORDIC.scala 454:32]
  wire [63:0] _fxxterm_T_31 = 64'sh0 - $signed(x_7); // @[VCORDIC.scala 454:45]
  wire [63:0] fxxterm_7 = $signed(y_7) < 64'sh0 ? $signed(_fxxterm_T_31) : $signed(x_7); // @[VCORDIC.scala 454:26]
  wire [63:0] _fxyterm_T_31 = 64'sh0 - $signed(y_7); // @[VCORDIC.scala 455:45]
  wire [63:0] fxyterm_7 = _fxxterm_T_28 ? $signed(_fxyterm_T_31) : $signed(y_7); // @[VCORDIC.scala 455:26]
  wire [63:0] _fxthetaterm_T_23 = 64'h0 - 64'h1fffd56; // @[VCORDIC.scala 456:49]
  wire [56:0] _GEN_12 = fxyterm_7[63:7]; // @[VCORDIC.scala 458:37]
  wire [63:0] _x_8_T = {{7{_GEN_12[56]}},_GEN_12}; // @[VCORDIC.scala 458:37]
  wire [63:0] x_8 = $signed(x_7) + $signed(_x_8_T); // @[VCORDIC.scala 458:26]
  wire [56:0] _GEN_13 = fxxterm_7[63:7]; // @[VCORDIC.scala 459:37]
  wire [63:0] _y_8_T = {{7{_GEN_13[56]}},_GEN_13}; // @[VCORDIC.scala 459:37]
  wire [63:0] y_8 = $signed(y_7) - $signed(_y_8_T); // @[VCORDIC.scala 459:26]
  wire [63:0] _z_8_T = _fxxterm_T_28 ? _fxthetaterm_T_23 : 64'h1fffd56; // @[VCORDIC.scala 460:40]
  wire [63:0] z_8 = $signed(z_7) + $signed(_z_8_T); // @[VCORDIC.scala 460:26]
  wire  _fxxterm_T_32 = $signed(y_8) < 64'sh0; // @[VCORDIC.scala 454:32]
  wire [63:0] _fxxterm_T_35 = 64'sh0 - $signed(x_8); // @[VCORDIC.scala 454:45]
  wire [63:0] fxxterm_8 = $signed(y_8) < 64'sh0 ? $signed(_fxxterm_T_35) : $signed(x_8); // @[VCORDIC.scala 454:26]
  wire [63:0] _fxyterm_T_35 = 64'sh0 - $signed(y_8); // @[VCORDIC.scala 455:45]
  wire [63:0] fxyterm_8 = _fxxterm_T_32 ? $signed(_fxyterm_T_35) : $signed(y_8); // @[VCORDIC.scala 455:26]
  wire [63:0] _fxthetaterm_T_26 = 64'h0 - 64'hffffab; // @[VCORDIC.scala 456:49]
  wire [55:0] _GEN_14 = fxyterm_8[63:8]; // @[VCORDIC.scala 458:37]
  wire [63:0] _x_9_T = {{8{_GEN_14[55]}},_GEN_14}; // @[VCORDIC.scala 458:37]
  wire [63:0] x_9 = $signed(x_8) + $signed(_x_9_T); // @[VCORDIC.scala 458:26]
  wire [55:0] _GEN_15 = fxxterm_8[63:8]; // @[VCORDIC.scala 459:37]
  wire [63:0] _y_9_T = {{8{_GEN_15[55]}},_GEN_15}; // @[VCORDIC.scala 459:37]
  wire [63:0] y_9 = $signed(y_8) - $signed(_y_9_T); // @[VCORDIC.scala 459:26]
  wire [63:0] _z_9_T = _fxxterm_T_32 ? _fxthetaterm_T_26 : 64'hffffab; // @[VCORDIC.scala 460:40]
  wire [63:0] z_9 = $signed(z_8) + $signed(_z_9_T); // @[VCORDIC.scala 460:26]
  wire  _fxxterm_T_36 = $signed(y_9) < 64'sh0; // @[VCORDIC.scala 454:32]
  wire [63:0] _fxxterm_T_39 = 64'sh0 - $signed(x_9); // @[VCORDIC.scala 454:45]
  wire [63:0] fxxterm_9 = $signed(y_9) < 64'sh0 ? $signed(_fxxterm_T_39) : $signed(x_9); // @[VCORDIC.scala 454:26]
  wire [63:0] _fxyterm_T_39 = 64'sh0 - $signed(y_9); // @[VCORDIC.scala 455:45]
  wire [63:0] fxyterm_9 = _fxxterm_T_36 ? $signed(_fxyterm_T_39) : $signed(y_9); // @[VCORDIC.scala 455:26]
  wire [63:0] _fxthetaterm_T_29 = 64'h0 - 64'h7ffff5; // @[VCORDIC.scala 456:49]
  wire [54:0] _GEN_16 = fxyterm_9[63:9]; // @[VCORDIC.scala 458:37]
  wire [63:0] _x_10_T = {{9{_GEN_16[54]}},_GEN_16}; // @[VCORDIC.scala 458:37]
  wire [63:0] x_10 = $signed(x_9) + $signed(_x_10_T); // @[VCORDIC.scala 458:26]
  wire [54:0] _GEN_17 = fxxterm_9[63:9]; // @[VCORDIC.scala 459:37]
  wire [63:0] _y_10_T = {{9{_GEN_17[54]}},_GEN_17}; // @[VCORDIC.scala 459:37]
  wire [63:0] y_10 = $signed(y_9) - $signed(_y_10_T); // @[VCORDIC.scala 459:26]
  wire [63:0] _z_10_T = _fxxterm_T_36 ? _fxthetaterm_T_29 : 64'h7ffff5; // @[VCORDIC.scala 460:40]
  wire [63:0] z_10 = $signed(z_9) + $signed(_z_10_T); // @[VCORDIC.scala 460:26]
  wire  _fxxterm_T_40 = $signed(y_10) < 64'sh0; // @[VCORDIC.scala 454:32]
  wire [63:0] _fxxterm_T_43 = 64'sh0 - $signed(x_10); // @[VCORDIC.scala 454:45]
  wire [63:0] fxxterm_10 = $signed(y_10) < 64'sh0 ? $signed(_fxxterm_T_43) : $signed(x_10); // @[VCORDIC.scala 454:26]
  wire [63:0] _fxyterm_T_43 = 64'sh0 - $signed(y_10); // @[VCORDIC.scala 455:45]
  wire [63:0] fxyterm_10 = _fxxterm_T_40 ? $signed(_fxyterm_T_43) : $signed(y_10); // @[VCORDIC.scala 455:26]
  wire [63:0] _fxthetaterm_T_32 = 64'h0 - 64'h3ffffe; // @[VCORDIC.scala 456:49]
  wire [53:0] _GEN_18 = fxyterm_10[63:10]; // @[VCORDIC.scala 458:37]
  wire [63:0] _x_11_T = {{10{_GEN_18[53]}},_GEN_18}; // @[VCORDIC.scala 458:37]
  wire [63:0] x_11 = $signed(x_10) + $signed(_x_11_T); // @[VCORDIC.scala 458:26]
  wire [53:0] _GEN_19 = fxxterm_10[63:10]; // @[VCORDIC.scala 459:37]
  wire [63:0] _y_11_T = {{10{_GEN_19[53]}},_GEN_19}; // @[VCORDIC.scala 459:37]
  wire [63:0] y_11 = $signed(y_10) - $signed(_y_11_T); // @[VCORDIC.scala 459:26]
  wire [63:0] _z_11_T = _fxxterm_T_40 ? _fxthetaterm_T_32 : 64'h3ffffe; // @[VCORDIC.scala 460:40]
  wire [63:0] z_11 = $signed(z_10) + $signed(_z_11_T); // @[VCORDIC.scala 460:26]
  wire  _fxxterm_T_44 = $signed(y_11) < 64'sh0; // @[VCORDIC.scala 454:32]
  wire [63:0] _fxxterm_T_47 = 64'sh0 - $signed(x_11); // @[VCORDIC.scala 454:45]
  wire [63:0] fxxterm_11 = $signed(y_11) < 64'sh0 ? $signed(_fxxterm_T_47) : $signed(x_11); // @[VCORDIC.scala 454:26]
  wire [63:0] _fxyterm_T_47 = 64'sh0 - $signed(y_11); // @[VCORDIC.scala 455:45]
  wire [63:0] fxyterm_11 = _fxxterm_T_44 ? $signed(_fxyterm_T_47) : $signed(y_11); // @[VCORDIC.scala 455:26]
  wire [63:0] _fxthetaterm_T_35 = 64'h0 - 64'h1fffff; // @[VCORDIC.scala 456:49]
  wire [52:0] _GEN_20 = fxyterm_11[63:11]; // @[VCORDIC.scala 458:37]
  wire [63:0] _x_12_T = {{11{_GEN_20[52]}},_GEN_20}; // @[VCORDIC.scala 458:37]
  wire [63:0] x_12 = $signed(x_11) + $signed(_x_12_T); // @[VCORDIC.scala 458:26]
  wire [52:0] _GEN_21 = fxxterm_11[63:11]; // @[VCORDIC.scala 459:37]
  wire [63:0] _y_12_T = {{11{_GEN_21[52]}},_GEN_21}; // @[VCORDIC.scala 459:37]
  wire [63:0] y_12 = $signed(y_11) - $signed(_y_12_T); // @[VCORDIC.scala 459:26]
  wire [63:0] _z_12_T = _fxxterm_T_44 ? _fxthetaterm_T_35 : 64'h1fffff; // @[VCORDIC.scala 460:40]
  wire [63:0] z_12 = $signed(z_11) + $signed(_z_12_T); // @[VCORDIC.scala 460:26]
  wire  _fxxterm_T_48 = $signed(y_12) < 64'sh0; // @[VCORDIC.scala 454:32]
  wire [63:0] _fxxterm_T_51 = 64'sh0 - $signed(x_12); // @[VCORDIC.scala 454:45]
  wire [63:0] fxxterm_12 = $signed(y_12) < 64'sh0 ? $signed(_fxxterm_T_51) : $signed(x_12); // @[VCORDIC.scala 454:26]
  wire [63:0] _fxyterm_T_51 = 64'sh0 - $signed(y_12); // @[VCORDIC.scala 455:45]
  wire [63:0] fxyterm_12 = _fxxterm_T_48 ? $signed(_fxyterm_T_51) : $signed(y_12); // @[VCORDIC.scala 455:26]
  wire [63:0] _fxthetaterm_T_38 = 64'h0 - 64'h100000; // @[VCORDIC.scala 456:49]
  wire [51:0] _GEN_22 = fxyterm_12[63:12]; // @[VCORDIC.scala 458:37]
  wire [63:0] _x_13_T = {{12{_GEN_22[51]}},_GEN_22}; // @[VCORDIC.scala 458:37]
  wire [63:0] x_13 = $signed(x_12) + $signed(_x_13_T); // @[VCORDIC.scala 458:26]
  wire [51:0] _GEN_23 = fxxterm_12[63:12]; // @[VCORDIC.scala 459:37]
  wire [63:0] _y_13_T = {{12{_GEN_23[51]}},_GEN_23}; // @[VCORDIC.scala 459:37]
  wire [63:0] y_13 = $signed(y_12) - $signed(_y_13_T); // @[VCORDIC.scala 459:26]
  wire [63:0] _z_13_T = _fxxterm_T_48 ? _fxthetaterm_T_38 : 64'h100000; // @[VCORDIC.scala 460:40]
  wire [63:0] z_13 = $signed(z_12) + $signed(_z_13_T); // @[VCORDIC.scala 460:26]
  wire  _fxxterm_T_52 = $signed(y_13) < 64'sh0; // @[VCORDIC.scala 454:32]
  wire [63:0] _fxxterm_T_55 = 64'sh0 - $signed(x_13); // @[VCORDIC.scala 454:45]
  wire [63:0] fxxterm_13 = $signed(y_13) < 64'sh0 ? $signed(_fxxterm_T_55) : $signed(x_13); // @[VCORDIC.scala 454:26]
  wire [63:0] _fxyterm_T_55 = 64'sh0 - $signed(y_13); // @[VCORDIC.scala 455:45]
  wire [63:0] fxyterm_13 = _fxxterm_T_52 ? $signed(_fxyterm_T_55) : $signed(y_13); // @[VCORDIC.scala 455:26]
  wire [63:0] _fxthetaterm_T_41 = 64'h0 - 64'h80000; // @[VCORDIC.scala 456:49]
  wire [50:0] _GEN_24 = fxyterm_13[63:13]; // @[VCORDIC.scala 458:37]
  wire [63:0] _x_14_T = {{13{_GEN_24[50]}},_GEN_24}; // @[VCORDIC.scala 458:37]
  wire [63:0] x_14 = $signed(x_13) + $signed(_x_14_T); // @[VCORDIC.scala 458:26]
  wire [50:0] _GEN_25 = fxxterm_13[63:13]; // @[VCORDIC.scala 459:37]
  wire [63:0] _y_14_T = {{13{_GEN_25[50]}},_GEN_25}; // @[VCORDIC.scala 459:37]
  wire [63:0] y_14 = $signed(y_13) - $signed(_y_14_T); // @[VCORDIC.scala 459:26]
  wire [63:0] _z_14_T = _fxxterm_T_52 ? _fxthetaterm_T_41 : 64'h80000; // @[VCORDIC.scala 460:40]
  wire [63:0] z_14 = $signed(z_13) + $signed(_z_14_T); // @[VCORDIC.scala 460:26]
  wire  _fxxterm_T_56 = $signed(y_14) < 64'sh0; // @[VCORDIC.scala 454:32]
  wire [63:0] _fxxterm_T_59 = 64'sh0 - $signed(x_14); // @[VCORDIC.scala 454:45]
  wire [63:0] fxxterm_14 = $signed(y_14) < 64'sh0 ? $signed(_fxxterm_T_59) : $signed(x_14); // @[VCORDIC.scala 454:26]
  wire [63:0] _fxyterm_T_59 = 64'sh0 - $signed(y_14); // @[VCORDIC.scala 455:45]
  wire [63:0] fxyterm_14 = _fxxterm_T_56 ? $signed(_fxyterm_T_59) : $signed(y_14); // @[VCORDIC.scala 455:26]
  wire [63:0] _fxthetaterm_T_44 = 64'h0 - 64'h40000; // @[VCORDIC.scala 456:49]
  wire [49:0] _GEN_26 = fxyterm_14[63:14]; // @[VCORDIC.scala 458:37]
  wire [63:0] _x_15_T = {{14{_GEN_26[49]}},_GEN_26}; // @[VCORDIC.scala 458:37]
  wire [63:0] x_15 = $signed(x_14) + $signed(_x_15_T); // @[VCORDIC.scala 458:26]
  wire [49:0] _GEN_27 = fxxterm_14[63:14]; // @[VCORDIC.scala 459:37]
  wire [63:0] _y_15_T = {{14{_GEN_27[49]}},_GEN_27}; // @[VCORDIC.scala 459:37]
  wire [63:0] y_15 = $signed(y_14) - $signed(_y_15_T); // @[VCORDIC.scala 459:26]
  wire [63:0] _z_15_T = _fxxterm_T_56 ? _fxthetaterm_T_44 : 64'h40000; // @[VCORDIC.scala 460:40]
  wire [63:0] z_15 = $signed(z_14) + $signed(_z_15_T); // @[VCORDIC.scala 460:26]
  wire  _fxxterm_T_60 = $signed(y_15) < 64'sh0; // @[VCORDIC.scala 454:32]
  wire [63:0] _fxxterm_T_63 = 64'sh0 - $signed(x_15); // @[VCORDIC.scala 454:45]
  wire [63:0] fxxterm_15 = $signed(y_15) < 64'sh0 ? $signed(_fxxterm_T_63) : $signed(x_15); // @[VCORDIC.scala 454:26]
  wire [63:0] _fxyterm_T_63 = 64'sh0 - $signed(y_15); // @[VCORDIC.scala 455:45]
  wire [63:0] fxyterm_15 = _fxxterm_T_60 ? $signed(_fxyterm_T_63) : $signed(y_15); // @[VCORDIC.scala 455:26]
  wire [63:0] _fxthetaterm_T_47 = 64'h0 - 64'h20000; // @[VCORDIC.scala 456:49]
  wire [48:0] _GEN_28 = fxyterm_15[63:15]; // @[VCORDIC.scala 458:37]
  wire [63:0] _x_16_T = {{15{_GEN_28[48]}},_GEN_28}; // @[VCORDIC.scala 458:37]
  wire [63:0] x_16 = $signed(x_15) + $signed(_x_16_T); // @[VCORDIC.scala 458:26]
  wire [48:0] _GEN_29 = fxxterm_15[63:15]; // @[VCORDIC.scala 459:37]
  wire [63:0] _y_16_T = {{15{_GEN_29[48]}},_GEN_29}; // @[VCORDIC.scala 459:37]
  wire [63:0] y_16 = $signed(y_15) - $signed(_y_16_T); // @[VCORDIC.scala 459:26]
  wire [63:0] _z_16_T = _fxxterm_T_60 ? _fxthetaterm_T_47 : 64'h20000; // @[VCORDIC.scala 460:40]
  wire [63:0] z_16 = $signed(z_15) + $signed(_z_16_T); // @[VCORDIC.scala 460:26]
  wire  _fxxterm_T_64 = $signed(y_16) < 64'sh0; // @[VCORDIC.scala 454:32]
  wire [63:0] _fxxterm_T_67 = 64'sh0 - $signed(x_16); // @[VCORDIC.scala 454:45]
  wire [63:0] fxxterm_16 = $signed(y_16) < 64'sh0 ? $signed(_fxxterm_T_67) : $signed(x_16); // @[VCORDIC.scala 454:26]
  wire [63:0] _fxyterm_T_67 = 64'sh0 - $signed(y_16); // @[VCORDIC.scala 455:45]
  wire [63:0] fxyterm_16 = _fxxterm_T_64 ? $signed(_fxyterm_T_67) : $signed(y_16); // @[VCORDIC.scala 455:26]
  wire [63:0] _fxthetaterm_T_50 = 64'h0 - 64'h10000; // @[VCORDIC.scala 456:49]
  wire [47:0] _GEN_30 = fxyterm_16[63:16]; // @[VCORDIC.scala 458:37]
  wire [63:0] _x_17_T = {{16{_GEN_30[47]}},_GEN_30}; // @[VCORDIC.scala 458:37]
  wire [63:0] x_17 = $signed(x_16) + $signed(_x_17_T); // @[VCORDIC.scala 458:26]
  wire [47:0] _GEN_31 = fxxterm_16[63:16]; // @[VCORDIC.scala 459:37]
  wire [63:0] _y_17_T = {{16{_GEN_31[47]}},_GEN_31}; // @[VCORDIC.scala 459:37]
  wire [63:0] y_17 = $signed(y_16) - $signed(_y_17_T); // @[VCORDIC.scala 459:26]
  wire [63:0] _z_17_T = _fxxterm_T_64 ? _fxthetaterm_T_50 : 64'h10000; // @[VCORDIC.scala 460:40]
  wire [63:0] z_17 = $signed(z_16) + $signed(_z_17_T); // @[VCORDIC.scala 460:26]
  wire  _fxxterm_T_68 = $signed(y_17) < 64'sh0; // @[VCORDIC.scala 454:32]
  wire [63:0] _fxxterm_T_71 = 64'sh0 - $signed(x_17); // @[VCORDIC.scala 454:45]
  wire [63:0] fxxterm_17 = $signed(y_17) < 64'sh0 ? $signed(_fxxterm_T_71) : $signed(x_17); // @[VCORDIC.scala 454:26]
  wire [63:0] _fxyterm_T_71 = 64'sh0 - $signed(y_17); // @[VCORDIC.scala 455:45]
  wire [63:0] fxyterm_17 = _fxxterm_T_68 ? $signed(_fxyterm_T_71) : $signed(y_17); // @[VCORDIC.scala 455:26]
  wire [63:0] _fxthetaterm_T_53 = 64'h0 - 64'h8000; // @[VCORDIC.scala 456:49]
  wire [46:0] _GEN_32 = fxyterm_17[63:17]; // @[VCORDIC.scala 458:37]
  wire [63:0] _x_18_T = {{17{_GEN_32[46]}},_GEN_32}; // @[VCORDIC.scala 458:37]
  wire [63:0] x_18 = $signed(x_17) + $signed(_x_18_T); // @[VCORDIC.scala 458:26]
  wire [46:0] _GEN_33 = fxxterm_17[63:17]; // @[VCORDIC.scala 459:37]
  wire [63:0] _y_18_T = {{17{_GEN_33[46]}},_GEN_33}; // @[VCORDIC.scala 459:37]
  wire [63:0] y_18 = $signed(y_17) - $signed(_y_18_T); // @[VCORDIC.scala 459:26]
  wire [63:0] _z_18_T = _fxxterm_T_68 ? _fxthetaterm_T_53 : 64'h8000; // @[VCORDIC.scala 460:40]
  wire [63:0] z_18 = $signed(z_17) + $signed(_z_18_T); // @[VCORDIC.scala 460:26]
  wire  _fxxterm_T_72 = $signed(y_18) < 64'sh0; // @[VCORDIC.scala 454:32]
  wire [63:0] _fxxterm_T_75 = 64'sh0 - $signed(x_18); // @[VCORDIC.scala 454:45]
  wire [63:0] fxxterm_18 = $signed(y_18) < 64'sh0 ? $signed(_fxxterm_T_75) : $signed(x_18); // @[VCORDIC.scala 454:26]
  wire [63:0] _fxyterm_T_75 = 64'sh0 - $signed(y_18); // @[VCORDIC.scala 455:45]
  wire [63:0] fxyterm_18 = _fxxterm_T_72 ? $signed(_fxyterm_T_75) : $signed(y_18); // @[VCORDIC.scala 455:26]
  wire [63:0] _fxthetaterm_T_56 = 64'h0 - 64'h4000; // @[VCORDIC.scala 456:49]
  wire [45:0] _GEN_34 = fxyterm_18[63:18]; // @[VCORDIC.scala 458:37]
  wire [63:0] _x_19_T = {{18{_GEN_34[45]}},_GEN_34}; // @[VCORDIC.scala 458:37]
  wire [63:0] x_19 = $signed(x_18) + $signed(_x_19_T); // @[VCORDIC.scala 458:26]
  wire [45:0] _GEN_35 = fxxterm_18[63:18]; // @[VCORDIC.scala 459:37]
  wire [63:0] _y_19_T = {{18{_GEN_35[45]}},_GEN_35}; // @[VCORDIC.scala 459:37]
  wire [63:0] y_19 = $signed(y_18) - $signed(_y_19_T); // @[VCORDIC.scala 459:26]
  wire [63:0] _z_19_T = _fxxterm_T_72 ? _fxthetaterm_T_56 : 64'h4000; // @[VCORDIC.scala 460:40]
  wire [63:0] z_19 = $signed(z_18) + $signed(_z_19_T); // @[VCORDIC.scala 460:26]
  wire  _fxxterm_T_76 = $signed(y_19) < 64'sh0; // @[VCORDIC.scala 454:32]
  wire [63:0] _fxxterm_T_79 = 64'sh0 - $signed(x_19); // @[VCORDIC.scala 454:45]
  wire [63:0] fxxterm_19 = $signed(y_19) < 64'sh0 ? $signed(_fxxterm_T_79) : $signed(x_19); // @[VCORDIC.scala 454:26]
  wire [63:0] _fxyterm_T_79 = 64'sh0 - $signed(y_19); // @[VCORDIC.scala 455:45]
  wire [63:0] fxyterm_19 = _fxxterm_T_76 ? $signed(_fxyterm_T_79) : $signed(y_19); // @[VCORDIC.scala 455:26]
  wire [63:0] _fxthetaterm_T_59 = 64'h0 - 64'h2000; // @[VCORDIC.scala 456:49]
  wire [44:0] _GEN_36 = fxyterm_19[63:19]; // @[VCORDIC.scala 458:37]
  wire [63:0] _x_20_T = {{19{_GEN_36[44]}},_GEN_36}; // @[VCORDIC.scala 458:37]
  wire [63:0] x_20 = $signed(x_19) + $signed(_x_20_T); // @[VCORDIC.scala 458:26]
  wire [44:0] _GEN_37 = fxxterm_19[63:19]; // @[VCORDIC.scala 459:37]
  wire [63:0] _y_20_T = {{19{_GEN_37[44]}},_GEN_37}; // @[VCORDIC.scala 459:37]
  wire [63:0] y_20 = $signed(y_19) - $signed(_y_20_T); // @[VCORDIC.scala 459:26]
  wire [63:0] _z_20_T = _fxxterm_T_76 ? _fxthetaterm_T_59 : 64'h2000; // @[VCORDIC.scala 460:40]
  wire [63:0] z_20 = $signed(z_19) + $signed(_z_20_T); // @[VCORDIC.scala 460:26]
  wire  _fxxterm_T_80 = $signed(y_20) < 64'sh0; // @[VCORDIC.scala 454:32]
  wire [63:0] _fxxterm_T_83 = 64'sh0 - $signed(x_20); // @[VCORDIC.scala 454:45]
  wire [63:0] fxxterm_20 = $signed(y_20) < 64'sh0 ? $signed(_fxxterm_T_83) : $signed(x_20); // @[VCORDIC.scala 454:26]
  wire [63:0] _fxyterm_T_83 = 64'sh0 - $signed(y_20); // @[VCORDIC.scala 455:45]
  wire [63:0] fxyterm_20 = _fxxterm_T_80 ? $signed(_fxyterm_T_83) : $signed(y_20); // @[VCORDIC.scala 455:26]
  wire [63:0] _fxthetaterm_T_62 = 64'h0 - 64'h1000; // @[VCORDIC.scala 456:49]
  wire [43:0] _GEN_38 = fxyterm_20[63:20]; // @[VCORDIC.scala 458:37]
  wire [63:0] _x_21_T = {{20{_GEN_38[43]}},_GEN_38}; // @[VCORDIC.scala 458:37]
  wire [63:0] x_21 = $signed(x_20) + $signed(_x_21_T); // @[VCORDIC.scala 458:26]
  wire [43:0] _GEN_39 = fxxterm_20[63:20]; // @[VCORDIC.scala 459:37]
  wire [63:0] _y_21_T = {{20{_GEN_39[43]}},_GEN_39}; // @[VCORDIC.scala 459:37]
  wire [63:0] y_21 = $signed(y_20) - $signed(_y_21_T); // @[VCORDIC.scala 459:26]
  wire [63:0] _z_21_T = _fxxterm_T_80 ? _fxthetaterm_T_62 : 64'h1000; // @[VCORDIC.scala 460:40]
  wire [63:0] z_21 = $signed(z_20) + $signed(_z_21_T); // @[VCORDIC.scala 460:26]
  wire  _fxxterm_T_84 = $signed(y_21) < 64'sh0; // @[VCORDIC.scala 454:32]
  wire [63:0] _fxxterm_T_87 = 64'sh0 - $signed(x_21); // @[VCORDIC.scala 454:45]
  wire [63:0] fxxterm_21 = $signed(y_21) < 64'sh0 ? $signed(_fxxterm_T_87) : $signed(x_21); // @[VCORDIC.scala 454:26]
  wire [63:0] _fxyterm_T_87 = 64'sh0 - $signed(y_21); // @[VCORDIC.scala 455:45]
  wire [63:0] fxyterm_21 = _fxxterm_T_84 ? $signed(_fxyterm_T_87) : $signed(y_21); // @[VCORDIC.scala 455:26]
  wire [63:0] _fxthetaterm_T_65 = 64'h0 - 64'h800; // @[VCORDIC.scala 456:49]
  wire [42:0] _GEN_40 = fxyterm_21[63:21]; // @[VCORDIC.scala 458:37]
  wire [63:0] _x_22_T = {{21{_GEN_40[42]}},_GEN_40}; // @[VCORDIC.scala 458:37]
  wire [63:0] x_22 = $signed(x_21) + $signed(_x_22_T); // @[VCORDIC.scala 458:26]
  wire [42:0] _GEN_41 = fxxterm_21[63:21]; // @[VCORDIC.scala 459:37]
  wire [63:0] _y_22_T = {{21{_GEN_41[42]}},_GEN_41}; // @[VCORDIC.scala 459:37]
  wire [63:0] y_22 = $signed(y_21) - $signed(_y_22_T); // @[VCORDIC.scala 459:26]
  wire [63:0] _z_22_T = _fxxterm_T_84 ? _fxthetaterm_T_65 : 64'h800; // @[VCORDIC.scala 460:40]
  wire [63:0] z_22 = $signed(z_21) + $signed(_z_22_T); // @[VCORDIC.scala 460:26]
  wire  _fxxterm_T_88 = $signed(y_22) < 64'sh0; // @[VCORDIC.scala 454:32]
  wire [63:0] _fxxterm_T_91 = 64'sh0 - $signed(x_22); // @[VCORDIC.scala 454:45]
  wire [63:0] fxxterm_22 = $signed(y_22) < 64'sh0 ? $signed(_fxxterm_T_91) : $signed(x_22); // @[VCORDIC.scala 454:26]
  wire [63:0] _fxyterm_T_91 = 64'sh0 - $signed(y_22); // @[VCORDIC.scala 455:45]
  wire [63:0] fxyterm_22 = _fxxterm_T_88 ? $signed(_fxyterm_T_91) : $signed(y_22); // @[VCORDIC.scala 455:26]
  wire [63:0] _fxthetaterm_T_68 = 64'h0 - 64'h400; // @[VCORDIC.scala 456:49]
  wire [41:0] _GEN_42 = fxyterm_22[63:22]; // @[VCORDIC.scala 458:37]
  wire [63:0] _x_23_T = {{22{_GEN_42[41]}},_GEN_42}; // @[VCORDIC.scala 458:37]
  wire [63:0] x_23 = $signed(x_22) + $signed(_x_23_T); // @[VCORDIC.scala 458:26]
  wire [41:0] _GEN_43 = fxxterm_22[63:22]; // @[VCORDIC.scala 459:37]
  wire [63:0] _y_23_T = {{22{_GEN_43[41]}},_GEN_43}; // @[VCORDIC.scala 459:37]
  wire [63:0] y_23 = $signed(y_22) - $signed(_y_23_T); // @[VCORDIC.scala 459:26]
  wire [63:0] _z_23_T = _fxxterm_T_88 ? _fxthetaterm_T_68 : 64'h400; // @[VCORDIC.scala 460:40]
  wire [63:0] z_23 = $signed(z_22) + $signed(_z_23_T); // @[VCORDIC.scala 460:26]
  wire  _fxxterm_T_92 = $signed(y_23) < 64'sh0; // @[VCORDIC.scala 454:32]
  wire [63:0] _fxxterm_T_95 = 64'sh0 - $signed(x_23); // @[VCORDIC.scala 454:45]
  wire [63:0] fxxterm_23 = $signed(y_23) < 64'sh0 ? $signed(_fxxterm_T_95) : $signed(x_23); // @[VCORDIC.scala 454:26]
  wire [63:0] _fxyterm_T_95 = 64'sh0 - $signed(y_23); // @[VCORDIC.scala 455:45]
  wire [63:0] fxyterm_23 = _fxxterm_T_92 ? $signed(_fxyterm_T_95) : $signed(y_23); // @[VCORDIC.scala 455:26]
  wire [63:0] _fxthetaterm_T_71 = 64'h0 - 64'h200; // @[VCORDIC.scala 456:49]
  wire [40:0] _GEN_44 = fxyterm_23[63:23]; // @[VCORDIC.scala 458:37]
  wire [63:0] _x_24_T = {{23{_GEN_44[40]}},_GEN_44}; // @[VCORDIC.scala 458:37]
  wire [63:0] x_24 = $signed(x_23) + $signed(_x_24_T); // @[VCORDIC.scala 458:26]
  wire [40:0] _GEN_45 = fxxterm_23[63:23]; // @[VCORDIC.scala 459:37]
  wire [63:0] _y_24_T = {{23{_GEN_45[40]}},_GEN_45}; // @[VCORDIC.scala 459:37]
  wire [63:0] y_24 = $signed(y_23) - $signed(_y_24_T); // @[VCORDIC.scala 459:26]
  wire [63:0] _z_24_T = _fxxterm_T_92 ? _fxthetaterm_T_71 : 64'h200; // @[VCORDIC.scala 460:40]
  wire [63:0] z_24 = $signed(z_23) + $signed(_z_24_T); // @[VCORDIC.scala 460:26]
  wire  _fxxterm_T_96 = $signed(y_24) < 64'sh0; // @[VCORDIC.scala 454:32]
  wire [63:0] _fxxterm_T_99 = 64'sh0 - $signed(x_24); // @[VCORDIC.scala 454:45]
  wire [63:0] fxxterm_24 = $signed(y_24) < 64'sh0 ? $signed(_fxxterm_T_99) : $signed(x_24); // @[VCORDIC.scala 454:26]
  wire [63:0] _fxyterm_T_99 = 64'sh0 - $signed(y_24); // @[VCORDIC.scala 455:45]
  wire [63:0] fxyterm_24 = _fxxterm_T_96 ? $signed(_fxyterm_T_99) : $signed(y_24); // @[VCORDIC.scala 455:26]
  wire [63:0] _fxthetaterm_T_74 = 64'h0 - 64'h100; // @[VCORDIC.scala 456:49]
  wire [39:0] _GEN_46 = fxyterm_24[63:24]; // @[VCORDIC.scala 458:37]
  wire [63:0] _x_25_T = {{24{_GEN_46[39]}},_GEN_46}; // @[VCORDIC.scala 458:37]
  wire [63:0] x_25 = $signed(x_24) + $signed(_x_25_T); // @[VCORDIC.scala 458:26]
  wire [39:0] _GEN_47 = fxxterm_24[63:24]; // @[VCORDIC.scala 459:37]
  wire [63:0] _y_25_T = {{24{_GEN_47[39]}},_GEN_47}; // @[VCORDIC.scala 459:37]
  wire [63:0] y_25 = $signed(y_24) - $signed(_y_25_T); // @[VCORDIC.scala 459:26]
  wire [63:0] _z_25_T = _fxxterm_T_96 ? _fxthetaterm_T_74 : 64'h100; // @[VCORDIC.scala 460:40]
  wire [63:0] z_25 = $signed(z_24) + $signed(_z_25_T); // @[VCORDIC.scala 460:26]
  wire  _fxxterm_T_100 = $signed(y_25) < 64'sh0; // @[VCORDIC.scala 454:32]
  wire [63:0] _fxxterm_T_103 = 64'sh0 - $signed(x_25); // @[VCORDIC.scala 454:45]
  wire [63:0] fxxterm_25 = $signed(y_25) < 64'sh0 ? $signed(_fxxterm_T_103) : $signed(x_25); // @[VCORDIC.scala 454:26]
  wire [63:0] _fxyterm_T_103 = 64'sh0 - $signed(y_25); // @[VCORDIC.scala 455:45]
  wire [63:0] fxyterm_25 = _fxxterm_T_100 ? $signed(_fxyterm_T_103) : $signed(y_25); // @[VCORDIC.scala 455:26]
  wire [63:0] _fxthetaterm_T_77 = 64'h0 - 64'h80; // @[VCORDIC.scala 456:49]
  wire [38:0] _GEN_48 = fxyterm_25[63:25]; // @[VCORDIC.scala 458:37]
  wire [63:0] _x_26_T = {{25{_GEN_48[38]}},_GEN_48}; // @[VCORDIC.scala 458:37]
  wire [63:0] x_26 = $signed(x_25) + $signed(_x_26_T); // @[VCORDIC.scala 458:26]
  wire [38:0] _GEN_49 = fxxterm_25[63:25]; // @[VCORDIC.scala 459:37]
  wire [63:0] _y_26_T = {{25{_GEN_49[38]}},_GEN_49}; // @[VCORDIC.scala 459:37]
  wire [63:0] y_26 = $signed(y_25) - $signed(_y_26_T); // @[VCORDIC.scala 459:26]
  wire [63:0] _z_26_T = _fxxterm_T_100 ? _fxthetaterm_T_77 : 64'h80; // @[VCORDIC.scala 460:40]
  wire [63:0] z_26 = $signed(z_25) + $signed(_z_26_T); // @[VCORDIC.scala 460:26]
  wire  _fxxterm_T_104 = $signed(y_26) < 64'sh0; // @[VCORDIC.scala 454:32]
  wire [63:0] _fxxterm_T_107 = 64'sh0 - $signed(x_26); // @[VCORDIC.scala 454:45]
  wire [63:0] fxxterm_26 = $signed(y_26) < 64'sh0 ? $signed(_fxxterm_T_107) : $signed(x_26); // @[VCORDIC.scala 454:26]
  wire [63:0] _fxyterm_T_107 = 64'sh0 - $signed(y_26); // @[VCORDIC.scala 455:45]
  wire [63:0] fxyterm_26 = _fxxterm_T_104 ? $signed(_fxyterm_T_107) : $signed(y_26); // @[VCORDIC.scala 455:26]
  wire [63:0] _fxthetaterm_T_80 = 64'h0 - 64'h40; // @[VCORDIC.scala 456:49]
  wire [37:0] _GEN_50 = fxyterm_26[63:26]; // @[VCORDIC.scala 458:37]
  wire [63:0] _x_27_T = {{26{_GEN_50[37]}},_GEN_50}; // @[VCORDIC.scala 458:37]
  wire [63:0] x_27 = $signed(x_26) + $signed(_x_27_T); // @[VCORDIC.scala 458:26]
  wire [37:0] _GEN_51 = fxxterm_26[63:26]; // @[VCORDIC.scala 459:37]
  wire [63:0] _y_27_T = {{26{_GEN_51[37]}},_GEN_51}; // @[VCORDIC.scala 459:37]
  wire [63:0] y_27 = $signed(y_26) - $signed(_y_27_T); // @[VCORDIC.scala 459:26]
  wire [63:0] _z_27_T = _fxxterm_T_104 ? _fxthetaterm_T_80 : 64'h40; // @[VCORDIC.scala 460:40]
  wire [63:0] z_27 = $signed(z_26) + $signed(_z_27_T); // @[VCORDIC.scala 460:26]
  wire  _fxxterm_T_108 = $signed(y_27) < 64'sh0; // @[VCORDIC.scala 454:32]
  wire [63:0] _fxxterm_T_111 = 64'sh0 - $signed(x_27); // @[VCORDIC.scala 454:45]
  wire [63:0] fxxterm_27 = $signed(y_27) < 64'sh0 ? $signed(_fxxterm_T_111) : $signed(x_27); // @[VCORDIC.scala 454:26]
  wire [63:0] _fxyterm_T_111 = 64'sh0 - $signed(y_27); // @[VCORDIC.scala 455:45]
  wire [63:0] fxyterm_27 = _fxxterm_T_108 ? $signed(_fxyterm_T_111) : $signed(y_27); // @[VCORDIC.scala 455:26]
  wire [63:0] _fxthetaterm_T_83 = 64'h0 - 64'h20; // @[VCORDIC.scala 456:49]
  wire [36:0] _GEN_52 = fxyterm_27[63:27]; // @[VCORDIC.scala 458:37]
  wire [63:0] _x_28_T = {{27{_GEN_52[36]}},_GEN_52}; // @[VCORDIC.scala 458:37]
  wire [63:0] x_28 = $signed(x_27) + $signed(_x_28_T); // @[VCORDIC.scala 458:26]
  wire [36:0] _GEN_53 = fxxterm_27[63:27]; // @[VCORDIC.scala 459:37]
  wire [63:0] _y_28_T = {{27{_GEN_53[36]}},_GEN_53}; // @[VCORDIC.scala 459:37]
  wire [63:0] y_28 = $signed(y_27) - $signed(_y_28_T); // @[VCORDIC.scala 459:26]
  wire [63:0] _z_28_T = _fxxterm_T_108 ? _fxthetaterm_T_83 : 64'h20; // @[VCORDIC.scala 460:40]
  wire [63:0] z_28 = $signed(z_27) + $signed(_z_28_T); // @[VCORDIC.scala 460:26]
  wire  _fxxterm_T_112 = $signed(y_28) < 64'sh0; // @[VCORDIC.scala 438:32]
  wire [63:0] _fxxterm_T_115 = 64'sh0 - $signed(x_28); // @[VCORDIC.scala 438:45]
  wire [63:0] fxxterm_28 = $signed(y_28) < 64'sh0 ? $signed(_fxxterm_T_115) : $signed(x_28); // @[VCORDIC.scala 438:26]
  wire [63:0] _fxyterm_T_115 = 64'sh0 - $signed(y_28); // @[VCORDIC.scala 439:45]
  wire [63:0] fxyterm_28 = _fxxterm_T_112 ? $signed(_fxyterm_T_115) : $signed(y_28); // @[VCORDIC.scala 439:26]
  wire [63:0] _fxthetaterm_T_86 = 64'h0 - 64'h10; // @[VCORDIC.scala 440:49]
  wire [35:0] _GEN_54 = fxyterm_28[63:28]; // @[VCORDIC.scala 442:37]
  wire [63:0] _x_29_T = {{28{_GEN_54[35]}},_GEN_54}; // @[VCORDIC.scala 442:37]
  wire [63:0] x_29 = $signed(x_28) + $signed(_x_29_T); // @[VCORDIC.scala 442:26]
  wire [35:0] _GEN_55 = fxxterm_28[63:28]; // @[VCORDIC.scala 443:37]
  wire [63:0] _y_29_T = {{28{_GEN_55[35]}},_GEN_55}; // @[VCORDIC.scala 443:37]
  wire [63:0] y_29 = $signed(y_28) - $signed(_y_29_T); // @[VCORDIC.scala 443:26]
  wire [63:0] _z_29_T = _fxxterm_T_112 ? _fxthetaterm_T_86 : 64'h10; // @[VCORDIC.scala 444:40]
  wire [63:0] z_29 = $signed(z_28) + $signed(_z_29_T); // @[VCORDIC.scala 444:26]
  Float32ToFixed64 tofixedx0 ( // @[VCORDIC.scala 107:33]
    .io_in(tofixedx0_io_in),
    .io_out(tofixedx0_io_out)
  );
  Float32ToFixed64 tofixedy0 ( // @[VCORDIC.scala 108:33]
    .io_in(tofixedy0_io_in),
    .io_out(tofixedy0_io_out)
  );
  Float32ToFixed64 tofixedz0 ( // @[VCORDIC.scala 109:33]
    .io_in(tofixedz0_io_in),
    .io_out(tofixedz0_io_out)
  );
  Fixed64ToFloat32 tofloatxout ( // @[VCORDIC.scala 467:29]
    .io_in(tofloatxout_io_in),
    .io_out(tofloatxout_io_out)
  );
  Fixed64ToFloat32 tofloatyout ( // @[VCORDIC.scala 468:29]
    .io_in(tofloatyout_io_in),
    .io_out(tofloatyout_io_out)
  );
  Fixed64ToFloat32 tofloatzout ( // @[VCORDIC.scala 469:29]
    .io_in(tofloatzout_io_in),
    .io_out(tofloatzout_io_out)
  );
  assign io_out_z = tofloatzout_io_out; // @[VCORDIC.scala 478:14]
  assign tofixedx0_io_in = 32'h3f800000; // @[VCORDIC.scala 111:19]
  assign tofixedy0_io_in = io_in_y0; // @[VCORDIC.scala 112:19]
  assign tofixedz0_io_in = 32'h0; // @[VCORDIC.scala 113:19]
  assign tofloatxout_io_in = xr_1; // @[VCORDIC.scala 472:32]
  assign tofloatyout_io_in = yr_1; // @[VCORDIC.scala 473:32]
  assign tofloatzout_io_in = zr_1; // @[VCORDIC.scala 474:32]
  always @(posedge clock) begin
    if (reset) begin // @[VCORDIC.scala 120:27]
      xr_0 <= 64'sh0; // @[VCORDIC.scala 120:27]
    end else begin
      xr_0 <= tofixedx0_io_out; // @[VCORDIC.scala 134:9]
    end
    if (reset) begin // @[VCORDIC.scala 120:27]
      xr_1 <= 64'sh0; // @[VCORDIC.scala 120:27]
    end else begin
      xr_1 <= x_29; // @[VCORDIC.scala 448:15]
    end
    if (reset) begin // @[VCORDIC.scala 121:27]
      yr_0 <= 64'sh0; // @[VCORDIC.scala 121:27]
    end else begin
      yr_0 <= tofixedy0_io_out; // @[VCORDIC.scala 135:9]
    end
    if (reset) begin // @[VCORDIC.scala 121:27]
      yr_1 <= 64'sh0; // @[VCORDIC.scala 121:27]
    end else begin
      yr_1 <= y_29; // @[VCORDIC.scala 449:15]
    end
    if (reset) begin // @[VCORDIC.scala 122:27]
      zr_0 <= 64'sh0; // @[VCORDIC.scala 122:27]
    end else begin
      zr_0 <= tofixedz0_io_out; // @[VCORDIC.scala 133:9]
    end
    if (reset) begin // @[VCORDIC.scala 122:27]
      zr_1 <= 64'sh0; // @[VCORDIC.scala 122:27]
    end else begin
      zr_1 <= z_29; // @[VCORDIC.scala 447:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  xr_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  xr_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  yr_0 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  yr_1 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  zr_0 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  zr_1 = _RAND_5[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
