module leadingOneDetector(
  input  [51:0] io_in,
  output [5:0]  io_out
);
  wire [1:0] _hotValue_T = io_in[1] ? 2'h2 : 2'h1; // @[Mux.scala 47:70]
  wire [1:0] _hotValue_T_1 = io_in[2] ? 2'h3 : _hotValue_T; // @[Mux.scala 47:70]
  wire [2:0] _hotValue_T_2 = io_in[3] ? 3'h4 : {{1'd0}, _hotValue_T_1}; // @[Mux.scala 47:70]
  wire [2:0] _hotValue_T_3 = io_in[4] ? 3'h5 : _hotValue_T_2; // @[Mux.scala 47:70]
  wire [2:0] _hotValue_T_4 = io_in[5] ? 3'h6 : _hotValue_T_3; // @[Mux.scala 47:70]
  wire [2:0] _hotValue_T_5 = io_in[6] ? 3'h7 : _hotValue_T_4; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_6 = io_in[7] ? 4'h8 : {{1'd0}, _hotValue_T_5}; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_7 = io_in[8] ? 4'h9 : _hotValue_T_6; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_8 = io_in[9] ? 4'ha : _hotValue_T_7; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_9 = io_in[10] ? 4'hb : _hotValue_T_8; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_10 = io_in[11] ? 4'hc : _hotValue_T_9; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_11 = io_in[12] ? 4'hd : _hotValue_T_10; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_12 = io_in[13] ? 4'he : _hotValue_T_11; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_13 = io_in[14] ? 4'hf : _hotValue_T_12; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_14 = io_in[15] ? 5'h10 : {{1'd0}, _hotValue_T_13}; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_15 = io_in[16] ? 5'h11 : _hotValue_T_14; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_16 = io_in[17] ? 5'h12 : _hotValue_T_15; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_17 = io_in[18] ? 5'h13 : _hotValue_T_16; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_18 = io_in[19] ? 5'h14 : _hotValue_T_17; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_19 = io_in[20] ? 5'h15 : _hotValue_T_18; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_20 = io_in[21] ? 5'h16 : _hotValue_T_19; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_21 = io_in[22] ? 5'h17 : _hotValue_T_20; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_22 = io_in[23] ? 5'h18 : _hotValue_T_21; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_23 = io_in[24] ? 5'h19 : _hotValue_T_22; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_24 = io_in[25] ? 5'h1a : _hotValue_T_23; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_25 = io_in[26] ? 5'h1b : _hotValue_T_24; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_26 = io_in[27] ? 5'h1c : _hotValue_T_25; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_27 = io_in[28] ? 5'h1d : _hotValue_T_26; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_28 = io_in[29] ? 5'h1e : _hotValue_T_27; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_29 = io_in[30] ? 5'h1f : _hotValue_T_28; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_30 = io_in[31] ? 6'h20 : {{1'd0}, _hotValue_T_29}; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_31 = io_in[32] ? 6'h21 : _hotValue_T_30; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_32 = io_in[33] ? 6'h22 : _hotValue_T_31; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_33 = io_in[34] ? 6'h23 : _hotValue_T_32; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_34 = io_in[35] ? 6'h24 : _hotValue_T_33; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_35 = io_in[36] ? 6'h25 : _hotValue_T_34; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_36 = io_in[37] ? 6'h26 : _hotValue_T_35; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_37 = io_in[38] ? 6'h27 : _hotValue_T_36; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_38 = io_in[39] ? 6'h28 : _hotValue_T_37; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_39 = io_in[40] ? 6'h29 : _hotValue_T_38; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_40 = io_in[41] ? 6'h2a : _hotValue_T_39; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_41 = io_in[42] ? 6'h2b : _hotValue_T_40; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_42 = io_in[43] ? 6'h2c : _hotValue_T_41; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_43 = io_in[44] ? 6'h2d : _hotValue_T_42; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_44 = io_in[45] ? 6'h2e : _hotValue_T_43; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_45 = io_in[46] ? 6'h2f : _hotValue_T_44; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_46 = io_in[47] ? 6'h30 : _hotValue_T_45; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_47 = io_in[48] ? 6'h31 : _hotValue_T_46; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_48 = io_in[49] ? 6'h32 : _hotValue_T_47; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_49 = io_in[50] ? 6'h33 : _hotValue_T_48; // @[Mux.scala 47:70]
  assign io_out = io_in[51] ? 6'h34 : _hotValue_T_49; // @[Mux.scala 47:70]
endmodule
