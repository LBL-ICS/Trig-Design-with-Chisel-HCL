module divider_BW106_v3(
  input          clock,
  input          reset,
  input  [105:0] io_in_a,
  output [105:0] io_out_s
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [127:0] _RAND_4;
  reg [127:0] _RAND_5;
  reg [127:0] _RAND_6;
  reg [127:0] _RAND_7;
  reg [127:0] _RAND_8;
  reg [127:0] _RAND_9;
  reg [127:0] _RAND_10;
  reg [127:0] _RAND_11;
  reg [127:0] _RAND_12;
  reg [127:0] _RAND_13;
  reg [127:0] _RAND_14;
  reg [127:0] _RAND_15;
  reg [127:0] _RAND_16;
  reg [127:0] _RAND_17;
  reg [127:0] _RAND_18;
  reg [127:0] _RAND_19;
  reg [127:0] _RAND_20;
  reg [127:0] _RAND_21;
  reg [127:0] _RAND_22;
  reg [127:0] _RAND_23;
  reg [127:0] _RAND_24;
  reg [127:0] _RAND_25;
  reg [127:0] _RAND_26;
  reg [127:0] _RAND_27;
  reg [127:0] _RAND_28;
  reg [127:0] _RAND_29;
  reg [127:0] _RAND_30;
  reg [127:0] _RAND_31;
  reg [127:0] _RAND_32;
  reg [127:0] _RAND_33;
  reg [127:0] _RAND_34;
  reg [127:0] _RAND_35;
  reg [127:0] _RAND_36;
  reg [127:0] _RAND_37;
  reg [127:0] _RAND_38;
  reg [127:0] _RAND_39;
  reg [127:0] _RAND_40;
  reg [127:0] _RAND_41;
  reg [127:0] _RAND_42;
  reg [127:0] _RAND_43;
  reg [127:0] _RAND_44;
  reg [127:0] _RAND_45;
  reg [127:0] _RAND_46;
  reg [127:0] _RAND_47;
  reg [127:0] _RAND_48;
  reg [127:0] _RAND_49;
  reg [127:0] _RAND_50;
  reg [127:0] _RAND_51;
  reg [127:0] _RAND_52;
  reg [127:0] _RAND_53;
  reg [127:0] _RAND_54;
  reg [127:0] _RAND_55;
  reg [127:0] _RAND_56;
  reg [127:0] _RAND_57;
  reg [127:0] _RAND_58;
  reg [127:0] _RAND_59;
  reg [127:0] _RAND_60;
  reg [127:0] _RAND_61;
  reg [127:0] _RAND_62;
  reg [127:0] _RAND_63;
  reg [127:0] _RAND_64;
  reg [127:0] _RAND_65;
  reg [127:0] _RAND_66;
  reg [127:0] _RAND_67;
  reg [127:0] _RAND_68;
  reg [127:0] _RAND_69;
  reg [127:0] _RAND_70;
  reg [127:0] _RAND_71;
  reg [127:0] _RAND_72;
  reg [127:0] _RAND_73;
  reg [127:0] _RAND_74;
  reg [127:0] _RAND_75;
  reg [127:0] _RAND_76;
  reg [127:0] _RAND_77;
  reg [127:0] _RAND_78;
  reg [127:0] _RAND_79;
  reg [127:0] _RAND_80;
  reg [127:0] _RAND_81;
  reg [127:0] _RAND_82;
  reg [127:0] _RAND_83;
  reg [127:0] _RAND_84;
  reg [127:0] _RAND_85;
  reg [127:0] _RAND_86;
  reg [127:0] _RAND_87;
  reg [127:0] _RAND_88;
  reg [127:0] _RAND_89;
  reg [127:0] _RAND_90;
  reg [127:0] _RAND_91;
  reg [127:0] _RAND_92;
  reg [127:0] _RAND_93;
  reg [127:0] _RAND_94;
  reg [127:0] _RAND_95;
  reg [127:0] _RAND_96;
  reg [127:0] _RAND_97;
  reg [127:0] _RAND_98;
  reg [127:0] _RAND_99;
  reg [127:0] _RAND_100;
  reg [127:0] _RAND_101;
  reg [127:0] _RAND_102;
  reg [127:0] _RAND_103;
  reg [127:0] _RAND_104;
  reg [127:0] _RAND_105;
  reg [127:0] _RAND_106;
  reg [127:0] _RAND_107;
  reg [127:0] _RAND_108;
  reg [127:0] _RAND_109;
  reg [127:0] _RAND_110;
  reg [127:0] _RAND_111;
  reg [127:0] _RAND_112;
  reg [127:0] _RAND_113;
  reg [127:0] _RAND_114;
  reg [127:0] _RAND_115;
  reg [127:0] _RAND_116;
  reg [127:0] _RAND_117;
  reg [127:0] _RAND_118;
  reg [127:0] _RAND_119;
  reg [127:0] _RAND_120;
  reg [127:0] _RAND_121;
  reg [127:0] _RAND_122;
  reg [127:0] _RAND_123;
  reg [127:0] _RAND_124;
  reg [127:0] _RAND_125;
  reg [127:0] _RAND_126;
  reg [127:0] _RAND_127;
  reg [127:0] _RAND_128;
  reg [127:0] _RAND_129;
  reg [127:0] _RAND_130;
  reg [127:0] _RAND_131;
  reg [127:0] _RAND_132;
  reg [127:0] _RAND_133;
  reg [127:0] _RAND_134;
  reg [127:0] _RAND_135;
  reg [127:0] _RAND_136;
  reg [127:0] _RAND_137;
  reg [127:0] _RAND_138;
  reg [127:0] _RAND_139;
  reg [127:0] _RAND_140;
  reg [127:0] _RAND_141;
  reg [127:0] _RAND_142;
  reg [127:0] _RAND_143;
  reg [127:0] _RAND_144;
  reg [127:0] _RAND_145;
  reg [127:0] _RAND_146;
  reg [127:0] _RAND_147;
  reg [127:0] _RAND_148;
  reg [127:0] _RAND_149;
  reg [127:0] _RAND_150;
  reg [127:0] _RAND_151;
  reg [127:0] _RAND_152;
  reg [127:0] _RAND_153;
  reg [127:0] _RAND_154;
  reg [127:0] _RAND_155;
`endif // RANDOMIZE_REG_INIT
  reg [105:0] a_aux_reg_r_0; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_1; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_2; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_3; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_4; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_5; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_6; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_7; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_8; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_9; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_10; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_11; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_12; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_13; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_14; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_15; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_16; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_17; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_18; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_19; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_20; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_21; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_22; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_23; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_24; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_25; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_26; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_27; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_28; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_29; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_30; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_31; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_32; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_33; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_34; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_35; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_36; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_37; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_38; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_39; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_40; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_41; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_42; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_43; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_44; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_45; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_46; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_47; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_48; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_49; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_50; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] a_aux_reg_r_51; // @[BinaryDesigns2.scala 171:30]
  reg [105:0] b_aux_reg_r_0; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_1; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_2; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_3; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_4; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_5; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_6; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_7; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_8; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_9; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_10; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_11; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_12; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_13; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_14; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_15; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_16; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_17; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_18; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_19; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_20; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_21; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_22; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_23; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_24; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_25; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_26; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_27; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_28; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_29; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_30; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_31; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_32; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_33; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_34; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_35; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_36; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_37; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_38; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_39; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_40; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_41; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_42; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_43; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_44; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_45; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_46; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_47; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_48; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_49; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_50; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] b_aux_reg_r_51; // @[BinaryDesigns2.scala 176:30]
  reg [105:0] result_reg_r_1; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_2; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_3; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_4; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_5; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_6; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_7; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_8; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_9; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_10; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_11; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_12; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_13; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_14; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_15; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_16; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_17; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_18; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_19; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_20; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_21; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_22; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_23; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_24; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_25; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_26; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_27; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_28; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_29; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_30; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_31; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_32; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_33; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_34; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_35; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_36; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_37; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_38; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_39; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_40; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_41; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_42; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_43; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_44; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_45; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_46; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_47; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_48; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_49; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_50; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_51; // @[BinaryDesigns2.scala 181:31]
  reg [105:0] result_reg_r_52; // @[BinaryDesigns2.scala 181:31]
  wire [208:0] _T_11240 = {b_aux_reg_r_0, 103'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [208:0] _GEN_1272 = {{103'd0}, a_aux_reg_r_0}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_1_103 = _GEN_1272 >= _T_11240; // @[BinaryDesigns2.scala 224:35]
  wire [105:0] result_reg_w_1 = {2'h0,wire_res_1_103,1'h0,3'h0,7'h0,13'h0,26'h0,53'h0}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_2_0 = result_reg_w_1[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_1 = result_reg_w_1[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_2 = result_reg_w_1[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_3 = result_reg_w_1[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_4 = result_reg_w_1[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_5 = result_reg_w_1[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_6 = result_reg_w_1[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_7 = result_reg_w_1[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_8 = result_reg_w_1[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_9 = result_reg_w_1[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_10 = result_reg_w_1[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_11 = result_reg_w_1[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_12 = result_reg_w_1[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_13 = result_reg_w_1[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_14 = result_reg_w_1[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_15 = result_reg_w_1[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_16 = result_reg_w_1[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_17 = result_reg_w_1[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_18 = result_reg_w_1[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_19 = result_reg_w_1[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_20 = result_reg_w_1[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_21 = result_reg_w_1[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_22 = result_reg_w_1[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_23 = result_reg_w_1[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_24 = result_reg_w_1[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_25 = result_reg_w_1[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_26 = result_reg_w_1[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_27 = result_reg_w_1[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_28 = result_reg_w_1[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_29 = result_reg_w_1[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_30 = result_reg_w_1[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_31 = result_reg_w_1[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_32 = result_reg_w_1[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_33 = result_reg_w_1[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_34 = result_reg_w_1[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_35 = result_reg_w_1[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_36 = result_reg_w_1[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_37 = result_reg_w_1[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_38 = result_reg_w_1[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_39 = result_reg_w_1[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_40 = result_reg_w_1[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_41 = result_reg_w_1[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_42 = result_reg_w_1[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_43 = result_reg_w_1[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_44 = result_reg_w_1[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_45 = result_reg_w_1[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_46 = result_reg_w_1[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_47 = result_reg_w_1[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_48 = result_reg_w_1[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_49 = result_reg_w_1[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_50 = result_reg_w_1[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_51 = result_reg_w_1[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_52 = result_reg_w_1[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_53 = result_reg_w_1[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_54 = result_reg_w_1[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_55 = result_reg_w_1[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_56 = result_reg_w_1[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_57 = result_reg_w_1[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_58 = result_reg_w_1[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_59 = result_reg_w_1[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_60 = result_reg_w_1[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_61 = result_reg_w_1[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_62 = result_reg_w_1[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_63 = result_reg_w_1[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_64 = result_reg_w_1[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_65 = result_reg_w_1[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_66 = result_reg_w_1[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_67 = result_reg_w_1[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_68 = result_reg_w_1[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_69 = result_reg_w_1[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_70 = result_reg_w_1[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_71 = result_reg_w_1[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_72 = result_reg_w_1[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_73 = result_reg_w_1[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_74 = result_reg_w_1[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_75 = result_reg_w_1[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_76 = result_reg_w_1[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_77 = result_reg_w_1[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_78 = result_reg_w_1[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_79 = result_reg_w_1[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_80 = result_reg_w_1[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_81 = result_reg_w_1[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_82 = result_reg_w_1[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_83 = result_reg_w_1[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_84 = result_reg_w_1[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_85 = result_reg_w_1[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_86 = result_reg_w_1[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_87 = result_reg_w_1[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_88 = result_reg_w_1[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_89 = result_reg_w_1[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_90 = result_reg_w_1[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_91 = result_reg_w_1[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_92 = result_reg_w_1[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_93 = result_reg_w_1[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_94 = result_reg_w_1[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_95 = result_reg_w_1[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_96 = result_reg_w_1[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_97 = result_reg_w_1[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_98 = result_reg_w_1[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_99 = result_reg_w_1[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_100 = result_reg_w_1[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_101 = result_reg_w_1[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_103 = result_reg_w_1[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_104 = result_reg_w_1[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_2_105 = result_reg_w_1[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_0 = result_reg_r_1[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_1 = result_reg_r_1[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_2 = result_reg_r_1[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_3 = result_reg_r_1[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_4 = result_reg_r_1[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_5 = result_reg_r_1[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_6 = result_reg_r_1[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_7 = result_reg_r_1[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_8 = result_reg_r_1[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_9 = result_reg_r_1[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_10 = result_reg_r_1[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_11 = result_reg_r_1[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_12 = result_reg_r_1[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_13 = result_reg_r_1[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_14 = result_reg_r_1[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_15 = result_reg_r_1[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_16 = result_reg_r_1[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_17 = result_reg_r_1[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_18 = result_reg_r_1[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_19 = result_reg_r_1[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_20 = result_reg_r_1[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_21 = result_reg_r_1[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_22 = result_reg_r_1[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_23 = result_reg_r_1[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_24 = result_reg_r_1[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_25 = result_reg_r_1[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_26 = result_reg_r_1[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_27 = result_reg_r_1[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_28 = result_reg_r_1[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_29 = result_reg_r_1[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_30 = result_reg_r_1[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_31 = result_reg_r_1[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_32 = result_reg_r_1[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_33 = result_reg_r_1[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_34 = result_reg_r_1[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_35 = result_reg_r_1[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_36 = result_reg_r_1[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_37 = result_reg_r_1[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_38 = result_reg_r_1[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_39 = result_reg_r_1[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_40 = result_reg_r_1[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_41 = result_reg_r_1[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_42 = result_reg_r_1[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_43 = result_reg_r_1[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_44 = result_reg_r_1[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_45 = result_reg_r_1[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_46 = result_reg_r_1[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_47 = result_reg_r_1[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_48 = result_reg_r_1[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_49 = result_reg_r_1[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_50 = result_reg_r_1[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_51 = result_reg_r_1[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_52 = result_reg_r_1[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_53 = result_reg_r_1[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_54 = result_reg_r_1[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_55 = result_reg_r_1[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_56 = result_reg_r_1[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_57 = result_reg_r_1[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_58 = result_reg_r_1[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_59 = result_reg_r_1[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_60 = result_reg_r_1[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_61 = result_reg_r_1[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_62 = result_reg_r_1[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_63 = result_reg_r_1[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_64 = result_reg_r_1[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_65 = result_reg_r_1[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_66 = result_reg_r_1[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_67 = result_reg_r_1[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_68 = result_reg_r_1[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_69 = result_reg_r_1[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_70 = result_reg_r_1[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_71 = result_reg_r_1[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_72 = result_reg_r_1[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_73 = result_reg_r_1[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_74 = result_reg_r_1[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_75 = result_reg_r_1[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_76 = result_reg_r_1[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_77 = result_reg_r_1[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_78 = result_reg_r_1[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_79 = result_reg_r_1[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_80 = result_reg_r_1[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_81 = result_reg_r_1[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_82 = result_reg_r_1[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_83 = result_reg_r_1[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_84 = result_reg_r_1[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_85 = result_reg_r_1[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_86 = result_reg_r_1[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_87 = result_reg_r_1[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_88 = result_reg_r_1[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_89 = result_reg_r_1[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_90 = result_reg_r_1[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_91 = result_reg_r_1[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_92 = result_reg_r_1[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_93 = result_reg_r_1[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_94 = result_reg_r_1[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_95 = result_reg_r_1[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_96 = result_reg_r_1[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_97 = result_reg_r_1[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_98 = result_reg_r_1[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_99 = result_reg_r_1[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_100 = result_reg_r_1[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_102 = result_reg_r_1[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_103 = result_reg_r_1[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_104 = result_reg_r_1[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_3_105 = result_reg_r_1[105]; // @[BinaryDesigns2.scala 192:62]
  wire [206:0] _T_11244 = {b_aux_reg_r_1, 101'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [206:0] _GEN_1273 = {{101'd0}, a_aux_reg_r_1}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_3_101 = _GEN_1273 >= _T_11244; // @[BinaryDesigns2.scala 224:35]
  wire [6:0] result_reg_w_2_hi_hi_hi_lo = {wire_res_3_98,wire_res_3_97,wire_res_3_96,wire_res_3_95,wire_res_3_94,
    wire_res_3_93,wire_res_3_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_2_hi_hi_lo_lo = {wire_res_3_84,wire_res_3_83,wire_res_3_82,wire_res_3_81,wire_res_3_80,
    wire_res_3_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_2_hi_hi_lo = {wire_res_3_91,wire_res_3_90,wire_res_3_89,wire_res_3_88,wire_res_3_87,
    wire_res_3_86,wire_res_3_85,result_reg_w_2_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_2_hi_lo_hi_lo = {wire_res_3_71,wire_res_3_70,wire_res_3_69,wire_res_3_68,wire_res_3_67,
    wire_res_3_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_2_hi_lo_lo_lo = {wire_res_3_58,wire_res_3_57,wire_res_3_56,wire_res_3_55,wire_res_3_54,
    wire_res_3_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_2_hi_lo_lo = {wire_res_3_65,wire_res_3_64,wire_res_3_63,wire_res_3_62,wire_res_3_61,
    wire_res_3_60,wire_res_3_59,result_reg_w_2_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_2_hi_lo = {wire_res_3_78,wire_res_3_77,wire_res_3_76,wire_res_3_75,wire_res_3_74,
    wire_res_3_73,wire_res_3_72,result_reg_w_2_hi_lo_hi_lo,result_reg_w_2_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_2_hi = {wire_res_3_105,wire_res_3_104,wire_res_3_103,wire_res_3_102,wire_res_3_101,
    wire_res_3_100,wire_res_3_99,result_reg_w_2_hi_hi_hi_lo,result_reg_w_2_hi_hi_lo,result_reg_w_2_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_2_lo_hi_hi_lo = {wire_res_3_45,wire_res_3_44,wire_res_3_43,wire_res_3_42,wire_res_3_41,
    wire_res_3_40,wire_res_3_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_2_lo_hi_lo_lo = {wire_res_3_31,wire_res_3_30,wire_res_3_29,wire_res_3_28,wire_res_3_27,
    wire_res_3_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_2_lo_hi_lo = {wire_res_3_38,wire_res_3_37,wire_res_3_36,wire_res_3_35,wire_res_3_34,
    wire_res_3_33,wire_res_3_32,result_reg_w_2_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_2_lo_lo_hi_lo = {wire_res_3_18,wire_res_3_17,wire_res_3_16,wire_res_3_15,wire_res_3_14,
    wire_res_3_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_2_lo_lo_lo_lo = {wire_res_3_5,wire_res_3_4,wire_res_3_3,wire_res_3_2,wire_res_3_1,wire_res_3_0
    }; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_2_lo_lo_lo = {wire_res_3_12,wire_res_3_11,wire_res_3_10,wire_res_3_9,wire_res_3_8,
    wire_res_3_7,wire_res_3_6,result_reg_w_2_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_2_lo_lo = {wire_res_3_25,wire_res_3_24,wire_res_3_23,wire_res_3_22,wire_res_3_21,
    wire_res_3_20,wire_res_3_19,result_reg_w_2_lo_lo_hi_lo,result_reg_w_2_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_2_lo = {wire_res_3_52,wire_res_3_51,wire_res_3_50,wire_res_3_49,wire_res_3_48,wire_res_3_47,
    wire_res_3_46,result_reg_w_2_lo_hi_hi_lo,result_reg_w_2_lo_hi_lo,result_reg_w_2_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_2 = {result_reg_w_2_hi,result_reg_w_2_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_4_0 = result_reg_w_2[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_1 = result_reg_w_2[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_2 = result_reg_w_2[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_3 = result_reg_w_2[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_4 = result_reg_w_2[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_5 = result_reg_w_2[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_6 = result_reg_w_2[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_7 = result_reg_w_2[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_8 = result_reg_w_2[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_9 = result_reg_w_2[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_10 = result_reg_w_2[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_11 = result_reg_w_2[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_12 = result_reg_w_2[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_13 = result_reg_w_2[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_14 = result_reg_w_2[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_15 = result_reg_w_2[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_16 = result_reg_w_2[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_17 = result_reg_w_2[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_18 = result_reg_w_2[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_19 = result_reg_w_2[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_20 = result_reg_w_2[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_21 = result_reg_w_2[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_22 = result_reg_w_2[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_23 = result_reg_w_2[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_24 = result_reg_w_2[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_25 = result_reg_w_2[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_26 = result_reg_w_2[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_27 = result_reg_w_2[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_28 = result_reg_w_2[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_29 = result_reg_w_2[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_30 = result_reg_w_2[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_31 = result_reg_w_2[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_32 = result_reg_w_2[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_33 = result_reg_w_2[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_34 = result_reg_w_2[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_35 = result_reg_w_2[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_36 = result_reg_w_2[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_37 = result_reg_w_2[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_38 = result_reg_w_2[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_39 = result_reg_w_2[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_40 = result_reg_w_2[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_41 = result_reg_w_2[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_42 = result_reg_w_2[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_43 = result_reg_w_2[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_44 = result_reg_w_2[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_45 = result_reg_w_2[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_46 = result_reg_w_2[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_47 = result_reg_w_2[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_48 = result_reg_w_2[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_49 = result_reg_w_2[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_50 = result_reg_w_2[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_51 = result_reg_w_2[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_52 = result_reg_w_2[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_53 = result_reg_w_2[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_54 = result_reg_w_2[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_55 = result_reg_w_2[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_56 = result_reg_w_2[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_57 = result_reg_w_2[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_58 = result_reg_w_2[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_59 = result_reg_w_2[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_60 = result_reg_w_2[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_61 = result_reg_w_2[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_62 = result_reg_w_2[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_63 = result_reg_w_2[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_64 = result_reg_w_2[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_65 = result_reg_w_2[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_66 = result_reg_w_2[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_67 = result_reg_w_2[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_68 = result_reg_w_2[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_69 = result_reg_w_2[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_70 = result_reg_w_2[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_71 = result_reg_w_2[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_72 = result_reg_w_2[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_73 = result_reg_w_2[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_74 = result_reg_w_2[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_75 = result_reg_w_2[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_76 = result_reg_w_2[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_77 = result_reg_w_2[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_78 = result_reg_w_2[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_79 = result_reg_w_2[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_80 = result_reg_w_2[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_81 = result_reg_w_2[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_82 = result_reg_w_2[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_83 = result_reg_w_2[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_84 = result_reg_w_2[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_85 = result_reg_w_2[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_86 = result_reg_w_2[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_87 = result_reg_w_2[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_88 = result_reg_w_2[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_89 = result_reg_w_2[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_90 = result_reg_w_2[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_91 = result_reg_w_2[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_92 = result_reg_w_2[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_93 = result_reg_w_2[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_94 = result_reg_w_2[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_95 = result_reg_w_2[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_96 = result_reg_w_2[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_97 = result_reg_w_2[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_98 = result_reg_w_2[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_99 = result_reg_w_2[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_101 = result_reg_w_2[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_102 = result_reg_w_2[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_103 = result_reg_w_2[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_104 = result_reg_w_2[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_4_105 = result_reg_w_2[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_0 = result_reg_r_2[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_1 = result_reg_r_2[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_2 = result_reg_r_2[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_3 = result_reg_r_2[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_4 = result_reg_r_2[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_5 = result_reg_r_2[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_6 = result_reg_r_2[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_7 = result_reg_r_2[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_8 = result_reg_r_2[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_9 = result_reg_r_2[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_10 = result_reg_r_2[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_11 = result_reg_r_2[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_12 = result_reg_r_2[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_13 = result_reg_r_2[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_14 = result_reg_r_2[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_15 = result_reg_r_2[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_16 = result_reg_r_2[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_17 = result_reg_r_2[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_18 = result_reg_r_2[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_19 = result_reg_r_2[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_20 = result_reg_r_2[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_21 = result_reg_r_2[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_22 = result_reg_r_2[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_23 = result_reg_r_2[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_24 = result_reg_r_2[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_25 = result_reg_r_2[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_26 = result_reg_r_2[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_27 = result_reg_r_2[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_28 = result_reg_r_2[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_29 = result_reg_r_2[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_30 = result_reg_r_2[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_31 = result_reg_r_2[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_32 = result_reg_r_2[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_33 = result_reg_r_2[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_34 = result_reg_r_2[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_35 = result_reg_r_2[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_36 = result_reg_r_2[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_37 = result_reg_r_2[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_38 = result_reg_r_2[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_39 = result_reg_r_2[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_40 = result_reg_r_2[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_41 = result_reg_r_2[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_42 = result_reg_r_2[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_43 = result_reg_r_2[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_44 = result_reg_r_2[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_45 = result_reg_r_2[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_46 = result_reg_r_2[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_47 = result_reg_r_2[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_48 = result_reg_r_2[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_49 = result_reg_r_2[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_50 = result_reg_r_2[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_51 = result_reg_r_2[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_52 = result_reg_r_2[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_53 = result_reg_r_2[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_54 = result_reg_r_2[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_55 = result_reg_r_2[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_56 = result_reg_r_2[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_57 = result_reg_r_2[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_58 = result_reg_r_2[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_59 = result_reg_r_2[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_60 = result_reg_r_2[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_61 = result_reg_r_2[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_62 = result_reg_r_2[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_63 = result_reg_r_2[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_64 = result_reg_r_2[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_65 = result_reg_r_2[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_66 = result_reg_r_2[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_67 = result_reg_r_2[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_68 = result_reg_r_2[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_69 = result_reg_r_2[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_70 = result_reg_r_2[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_71 = result_reg_r_2[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_72 = result_reg_r_2[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_73 = result_reg_r_2[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_74 = result_reg_r_2[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_75 = result_reg_r_2[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_76 = result_reg_r_2[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_77 = result_reg_r_2[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_78 = result_reg_r_2[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_79 = result_reg_r_2[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_80 = result_reg_r_2[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_81 = result_reg_r_2[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_82 = result_reg_r_2[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_83 = result_reg_r_2[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_84 = result_reg_r_2[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_85 = result_reg_r_2[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_86 = result_reg_r_2[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_87 = result_reg_r_2[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_88 = result_reg_r_2[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_89 = result_reg_r_2[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_90 = result_reg_r_2[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_91 = result_reg_r_2[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_92 = result_reg_r_2[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_93 = result_reg_r_2[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_94 = result_reg_r_2[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_95 = result_reg_r_2[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_96 = result_reg_r_2[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_97 = result_reg_r_2[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_98 = result_reg_r_2[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_100 = result_reg_r_2[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_101 = result_reg_r_2[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_102 = result_reg_r_2[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_103 = result_reg_r_2[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_104 = result_reg_r_2[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_5_105 = result_reg_r_2[105]; // @[BinaryDesigns2.scala 192:62]
  wire [204:0] _T_11248 = {b_aux_reg_r_2, 99'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [204:0] _GEN_1274 = {{99'd0}, a_aux_reg_r_2}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_5_99 = _GEN_1274 >= _T_11248; // @[BinaryDesigns2.scala 224:35]
  wire [6:0] result_reg_w_3_hi_hi_hi_lo = {wire_res_5_98,wire_res_5_97,wire_res_5_96,wire_res_5_95,wire_res_5_94,
    wire_res_5_93,wire_res_5_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_3_hi_hi_lo_lo = {wire_res_5_84,wire_res_5_83,wire_res_5_82,wire_res_5_81,wire_res_5_80,
    wire_res_5_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_3_hi_hi_lo = {wire_res_5_91,wire_res_5_90,wire_res_5_89,wire_res_5_88,wire_res_5_87,
    wire_res_5_86,wire_res_5_85,result_reg_w_3_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_3_hi_lo_hi_lo = {wire_res_5_71,wire_res_5_70,wire_res_5_69,wire_res_5_68,wire_res_5_67,
    wire_res_5_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_3_hi_lo_lo_lo = {wire_res_5_58,wire_res_5_57,wire_res_5_56,wire_res_5_55,wire_res_5_54,
    wire_res_5_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_3_hi_lo_lo = {wire_res_5_65,wire_res_5_64,wire_res_5_63,wire_res_5_62,wire_res_5_61,
    wire_res_5_60,wire_res_5_59,result_reg_w_3_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_3_hi_lo = {wire_res_5_78,wire_res_5_77,wire_res_5_76,wire_res_5_75,wire_res_5_74,
    wire_res_5_73,wire_res_5_72,result_reg_w_3_hi_lo_hi_lo,result_reg_w_3_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_3_hi = {wire_res_5_105,wire_res_5_104,wire_res_5_103,wire_res_5_102,wire_res_5_101,
    wire_res_5_100,wire_res_5_99,result_reg_w_3_hi_hi_hi_lo,result_reg_w_3_hi_hi_lo,result_reg_w_3_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_3_lo_hi_hi_lo = {wire_res_5_45,wire_res_5_44,wire_res_5_43,wire_res_5_42,wire_res_5_41,
    wire_res_5_40,wire_res_5_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_3_lo_hi_lo_lo = {wire_res_5_31,wire_res_5_30,wire_res_5_29,wire_res_5_28,wire_res_5_27,
    wire_res_5_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_3_lo_hi_lo = {wire_res_5_38,wire_res_5_37,wire_res_5_36,wire_res_5_35,wire_res_5_34,
    wire_res_5_33,wire_res_5_32,result_reg_w_3_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_3_lo_lo_hi_lo = {wire_res_5_18,wire_res_5_17,wire_res_5_16,wire_res_5_15,wire_res_5_14,
    wire_res_5_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_3_lo_lo_lo_lo = {wire_res_5_5,wire_res_5_4,wire_res_5_3,wire_res_5_2,wire_res_5_1,wire_res_5_0
    }; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_3_lo_lo_lo = {wire_res_5_12,wire_res_5_11,wire_res_5_10,wire_res_5_9,wire_res_5_8,
    wire_res_5_7,wire_res_5_6,result_reg_w_3_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_3_lo_lo = {wire_res_5_25,wire_res_5_24,wire_res_5_23,wire_res_5_22,wire_res_5_21,
    wire_res_5_20,wire_res_5_19,result_reg_w_3_lo_lo_hi_lo,result_reg_w_3_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_3_lo = {wire_res_5_52,wire_res_5_51,wire_res_5_50,wire_res_5_49,wire_res_5_48,wire_res_5_47,
    wire_res_5_46,result_reg_w_3_lo_hi_hi_lo,result_reg_w_3_lo_hi_lo,result_reg_w_3_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_3 = {result_reg_w_3_hi,result_reg_w_3_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_6_0 = result_reg_w_3[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_1 = result_reg_w_3[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_2 = result_reg_w_3[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_3 = result_reg_w_3[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_4 = result_reg_w_3[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_5 = result_reg_w_3[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_6 = result_reg_w_3[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_7 = result_reg_w_3[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_8 = result_reg_w_3[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_9 = result_reg_w_3[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_10 = result_reg_w_3[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_11 = result_reg_w_3[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_12 = result_reg_w_3[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_13 = result_reg_w_3[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_14 = result_reg_w_3[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_15 = result_reg_w_3[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_16 = result_reg_w_3[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_17 = result_reg_w_3[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_18 = result_reg_w_3[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_19 = result_reg_w_3[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_20 = result_reg_w_3[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_21 = result_reg_w_3[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_22 = result_reg_w_3[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_23 = result_reg_w_3[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_24 = result_reg_w_3[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_25 = result_reg_w_3[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_26 = result_reg_w_3[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_27 = result_reg_w_3[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_28 = result_reg_w_3[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_29 = result_reg_w_3[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_30 = result_reg_w_3[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_31 = result_reg_w_3[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_32 = result_reg_w_3[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_33 = result_reg_w_3[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_34 = result_reg_w_3[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_35 = result_reg_w_3[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_36 = result_reg_w_3[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_37 = result_reg_w_3[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_38 = result_reg_w_3[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_39 = result_reg_w_3[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_40 = result_reg_w_3[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_41 = result_reg_w_3[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_42 = result_reg_w_3[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_43 = result_reg_w_3[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_44 = result_reg_w_3[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_45 = result_reg_w_3[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_46 = result_reg_w_3[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_47 = result_reg_w_3[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_48 = result_reg_w_3[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_49 = result_reg_w_3[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_50 = result_reg_w_3[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_51 = result_reg_w_3[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_52 = result_reg_w_3[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_53 = result_reg_w_3[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_54 = result_reg_w_3[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_55 = result_reg_w_3[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_56 = result_reg_w_3[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_57 = result_reg_w_3[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_58 = result_reg_w_3[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_59 = result_reg_w_3[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_60 = result_reg_w_3[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_61 = result_reg_w_3[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_62 = result_reg_w_3[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_63 = result_reg_w_3[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_64 = result_reg_w_3[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_65 = result_reg_w_3[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_66 = result_reg_w_3[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_67 = result_reg_w_3[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_68 = result_reg_w_3[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_69 = result_reg_w_3[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_70 = result_reg_w_3[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_71 = result_reg_w_3[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_72 = result_reg_w_3[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_73 = result_reg_w_3[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_74 = result_reg_w_3[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_75 = result_reg_w_3[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_76 = result_reg_w_3[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_77 = result_reg_w_3[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_78 = result_reg_w_3[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_79 = result_reg_w_3[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_80 = result_reg_w_3[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_81 = result_reg_w_3[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_82 = result_reg_w_3[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_83 = result_reg_w_3[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_84 = result_reg_w_3[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_85 = result_reg_w_3[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_86 = result_reg_w_3[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_87 = result_reg_w_3[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_88 = result_reg_w_3[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_89 = result_reg_w_3[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_90 = result_reg_w_3[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_91 = result_reg_w_3[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_92 = result_reg_w_3[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_93 = result_reg_w_3[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_94 = result_reg_w_3[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_95 = result_reg_w_3[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_96 = result_reg_w_3[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_97 = result_reg_w_3[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_99 = result_reg_w_3[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_100 = result_reg_w_3[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_101 = result_reg_w_3[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_102 = result_reg_w_3[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_103 = result_reg_w_3[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_104 = result_reg_w_3[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_6_105 = result_reg_w_3[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_0 = result_reg_r_3[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_1 = result_reg_r_3[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_2 = result_reg_r_3[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_3 = result_reg_r_3[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_4 = result_reg_r_3[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_5 = result_reg_r_3[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_6 = result_reg_r_3[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_7 = result_reg_r_3[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_8 = result_reg_r_3[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_9 = result_reg_r_3[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_10 = result_reg_r_3[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_11 = result_reg_r_3[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_12 = result_reg_r_3[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_13 = result_reg_r_3[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_14 = result_reg_r_3[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_15 = result_reg_r_3[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_16 = result_reg_r_3[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_17 = result_reg_r_3[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_18 = result_reg_r_3[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_19 = result_reg_r_3[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_20 = result_reg_r_3[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_21 = result_reg_r_3[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_22 = result_reg_r_3[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_23 = result_reg_r_3[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_24 = result_reg_r_3[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_25 = result_reg_r_3[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_26 = result_reg_r_3[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_27 = result_reg_r_3[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_28 = result_reg_r_3[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_29 = result_reg_r_3[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_30 = result_reg_r_3[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_31 = result_reg_r_3[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_32 = result_reg_r_3[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_33 = result_reg_r_3[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_34 = result_reg_r_3[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_35 = result_reg_r_3[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_36 = result_reg_r_3[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_37 = result_reg_r_3[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_38 = result_reg_r_3[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_39 = result_reg_r_3[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_40 = result_reg_r_3[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_41 = result_reg_r_3[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_42 = result_reg_r_3[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_43 = result_reg_r_3[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_44 = result_reg_r_3[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_45 = result_reg_r_3[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_46 = result_reg_r_3[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_47 = result_reg_r_3[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_48 = result_reg_r_3[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_49 = result_reg_r_3[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_50 = result_reg_r_3[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_51 = result_reg_r_3[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_52 = result_reg_r_3[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_53 = result_reg_r_3[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_54 = result_reg_r_3[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_55 = result_reg_r_3[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_56 = result_reg_r_3[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_57 = result_reg_r_3[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_58 = result_reg_r_3[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_59 = result_reg_r_3[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_60 = result_reg_r_3[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_61 = result_reg_r_3[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_62 = result_reg_r_3[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_63 = result_reg_r_3[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_64 = result_reg_r_3[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_65 = result_reg_r_3[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_66 = result_reg_r_3[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_67 = result_reg_r_3[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_68 = result_reg_r_3[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_69 = result_reg_r_3[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_70 = result_reg_r_3[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_71 = result_reg_r_3[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_72 = result_reg_r_3[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_73 = result_reg_r_3[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_74 = result_reg_r_3[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_75 = result_reg_r_3[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_76 = result_reg_r_3[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_77 = result_reg_r_3[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_78 = result_reg_r_3[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_79 = result_reg_r_3[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_80 = result_reg_r_3[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_81 = result_reg_r_3[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_82 = result_reg_r_3[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_83 = result_reg_r_3[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_84 = result_reg_r_3[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_85 = result_reg_r_3[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_86 = result_reg_r_3[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_87 = result_reg_r_3[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_88 = result_reg_r_3[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_89 = result_reg_r_3[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_90 = result_reg_r_3[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_91 = result_reg_r_3[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_92 = result_reg_r_3[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_93 = result_reg_r_3[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_94 = result_reg_r_3[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_95 = result_reg_r_3[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_96 = result_reg_r_3[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_98 = result_reg_r_3[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_99 = result_reg_r_3[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_100 = result_reg_r_3[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_101 = result_reg_r_3[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_102 = result_reg_r_3[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_103 = result_reg_r_3[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_104 = result_reg_r_3[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_7_105 = result_reg_r_3[105]; // @[BinaryDesigns2.scala 192:62]
  wire [202:0] _T_11252 = {b_aux_reg_r_3, 97'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [202:0] _GEN_1275 = {{97'd0}, a_aux_reg_r_3}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_7_97 = _GEN_1275 >= _T_11252; // @[BinaryDesigns2.scala 224:35]
  wire [6:0] result_reg_w_4_hi_hi_hi_lo = {wire_res_7_98,wire_res_7_97,wire_res_7_96,wire_res_7_95,wire_res_7_94,
    wire_res_7_93,wire_res_7_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_4_hi_hi_lo_lo = {wire_res_7_84,wire_res_7_83,wire_res_7_82,wire_res_7_81,wire_res_7_80,
    wire_res_7_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_4_hi_hi_lo = {wire_res_7_91,wire_res_7_90,wire_res_7_89,wire_res_7_88,wire_res_7_87,
    wire_res_7_86,wire_res_7_85,result_reg_w_4_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_4_hi_lo_hi_lo = {wire_res_7_71,wire_res_7_70,wire_res_7_69,wire_res_7_68,wire_res_7_67,
    wire_res_7_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_4_hi_lo_lo_lo = {wire_res_7_58,wire_res_7_57,wire_res_7_56,wire_res_7_55,wire_res_7_54,
    wire_res_7_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_4_hi_lo_lo = {wire_res_7_65,wire_res_7_64,wire_res_7_63,wire_res_7_62,wire_res_7_61,
    wire_res_7_60,wire_res_7_59,result_reg_w_4_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_4_hi_lo = {wire_res_7_78,wire_res_7_77,wire_res_7_76,wire_res_7_75,wire_res_7_74,
    wire_res_7_73,wire_res_7_72,result_reg_w_4_hi_lo_hi_lo,result_reg_w_4_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_4_hi = {wire_res_7_105,wire_res_7_104,wire_res_7_103,wire_res_7_102,wire_res_7_101,
    wire_res_7_100,wire_res_7_99,result_reg_w_4_hi_hi_hi_lo,result_reg_w_4_hi_hi_lo,result_reg_w_4_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_4_lo_hi_hi_lo = {wire_res_7_45,wire_res_7_44,wire_res_7_43,wire_res_7_42,wire_res_7_41,
    wire_res_7_40,wire_res_7_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_4_lo_hi_lo_lo = {wire_res_7_31,wire_res_7_30,wire_res_7_29,wire_res_7_28,wire_res_7_27,
    wire_res_7_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_4_lo_hi_lo = {wire_res_7_38,wire_res_7_37,wire_res_7_36,wire_res_7_35,wire_res_7_34,
    wire_res_7_33,wire_res_7_32,result_reg_w_4_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_4_lo_lo_hi_lo = {wire_res_7_18,wire_res_7_17,wire_res_7_16,wire_res_7_15,wire_res_7_14,
    wire_res_7_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_4_lo_lo_lo_lo = {wire_res_7_5,wire_res_7_4,wire_res_7_3,wire_res_7_2,wire_res_7_1,wire_res_7_0
    }; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_4_lo_lo_lo = {wire_res_7_12,wire_res_7_11,wire_res_7_10,wire_res_7_9,wire_res_7_8,
    wire_res_7_7,wire_res_7_6,result_reg_w_4_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_4_lo_lo = {wire_res_7_25,wire_res_7_24,wire_res_7_23,wire_res_7_22,wire_res_7_21,
    wire_res_7_20,wire_res_7_19,result_reg_w_4_lo_lo_hi_lo,result_reg_w_4_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_4_lo = {wire_res_7_52,wire_res_7_51,wire_res_7_50,wire_res_7_49,wire_res_7_48,wire_res_7_47,
    wire_res_7_46,result_reg_w_4_lo_hi_hi_lo,result_reg_w_4_lo_hi_lo,result_reg_w_4_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_4 = {result_reg_w_4_hi,result_reg_w_4_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_8_0 = result_reg_w_4[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_1 = result_reg_w_4[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_2 = result_reg_w_4[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_3 = result_reg_w_4[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_4 = result_reg_w_4[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_5 = result_reg_w_4[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_6 = result_reg_w_4[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_7 = result_reg_w_4[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_8 = result_reg_w_4[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_9 = result_reg_w_4[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_10 = result_reg_w_4[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_11 = result_reg_w_4[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_12 = result_reg_w_4[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_13 = result_reg_w_4[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_14 = result_reg_w_4[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_15 = result_reg_w_4[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_16 = result_reg_w_4[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_17 = result_reg_w_4[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_18 = result_reg_w_4[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_19 = result_reg_w_4[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_20 = result_reg_w_4[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_21 = result_reg_w_4[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_22 = result_reg_w_4[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_23 = result_reg_w_4[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_24 = result_reg_w_4[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_25 = result_reg_w_4[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_26 = result_reg_w_4[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_27 = result_reg_w_4[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_28 = result_reg_w_4[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_29 = result_reg_w_4[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_30 = result_reg_w_4[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_31 = result_reg_w_4[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_32 = result_reg_w_4[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_33 = result_reg_w_4[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_34 = result_reg_w_4[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_35 = result_reg_w_4[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_36 = result_reg_w_4[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_37 = result_reg_w_4[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_38 = result_reg_w_4[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_39 = result_reg_w_4[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_40 = result_reg_w_4[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_41 = result_reg_w_4[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_42 = result_reg_w_4[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_43 = result_reg_w_4[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_44 = result_reg_w_4[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_45 = result_reg_w_4[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_46 = result_reg_w_4[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_47 = result_reg_w_4[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_48 = result_reg_w_4[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_49 = result_reg_w_4[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_50 = result_reg_w_4[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_51 = result_reg_w_4[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_52 = result_reg_w_4[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_53 = result_reg_w_4[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_54 = result_reg_w_4[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_55 = result_reg_w_4[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_56 = result_reg_w_4[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_57 = result_reg_w_4[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_58 = result_reg_w_4[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_59 = result_reg_w_4[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_60 = result_reg_w_4[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_61 = result_reg_w_4[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_62 = result_reg_w_4[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_63 = result_reg_w_4[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_64 = result_reg_w_4[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_65 = result_reg_w_4[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_66 = result_reg_w_4[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_67 = result_reg_w_4[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_68 = result_reg_w_4[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_69 = result_reg_w_4[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_70 = result_reg_w_4[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_71 = result_reg_w_4[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_72 = result_reg_w_4[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_73 = result_reg_w_4[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_74 = result_reg_w_4[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_75 = result_reg_w_4[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_76 = result_reg_w_4[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_77 = result_reg_w_4[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_78 = result_reg_w_4[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_79 = result_reg_w_4[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_80 = result_reg_w_4[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_81 = result_reg_w_4[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_82 = result_reg_w_4[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_83 = result_reg_w_4[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_84 = result_reg_w_4[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_85 = result_reg_w_4[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_86 = result_reg_w_4[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_87 = result_reg_w_4[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_88 = result_reg_w_4[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_89 = result_reg_w_4[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_90 = result_reg_w_4[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_91 = result_reg_w_4[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_92 = result_reg_w_4[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_93 = result_reg_w_4[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_94 = result_reg_w_4[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_95 = result_reg_w_4[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_97 = result_reg_w_4[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_98 = result_reg_w_4[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_99 = result_reg_w_4[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_100 = result_reg_w_4[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_101 = result_reg_w_4[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_102 = result_reg_w_4[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_103 = result_reg_w_4[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_104 = result_reg_w_4[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_8_105 = result_reg_w_4[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_0 = result_reg_r_4[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_1 = result_reg_r_4[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_2 = result_reg_r_4[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_3 = result_reg_r_4[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_4 = result_reg_r_4[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_5 = result_reg_r_4[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_6 = result_reg_r_4[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_7 = result_reg_r_4[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_8 = result_reg_r_4[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_9 = result_reg_r_4[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_10 = result_reg_r_4[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_11 = result_reg_r_4[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_12 = result_reg_r_4[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_13 = result_reg_r_4[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_14 = result_reg_r_4[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_15 = result_reg_r_4[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_16 = result_reg_r_4[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_17 = result_reg_r_4[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_18 = result_reg_r_4[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_19 = result_reg_r_4[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_20 = result_reg_r_4[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_21 = result_reg_r_4[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_22 = result_reg_r_4[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_23 = result_reg_r_4[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_24 = result_reg_r_4[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_25 = result_reg_r_4[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_26 = result_reg_r_4[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_27 = result_reg_r_4[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_28 = result_reg_r_4[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_29 = result_reg_r_4[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_30 = result_reg_r_4[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_31 = result_reg_r_4[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_32 = result_reg_r_4[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_33 = result_reg_r_4[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_34 = result_reg_r_4[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_35 = result_reg_r_4[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_36 = result_reg_r_4[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_37 = result_reg_r_4[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_38 = result_reg_r_4[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_39 = result_reg_r_4[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_40 = result_reg_r_4[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_41 = result_reg_r_4[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_42 = result_reg_r_4[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_43 = result_reg_r_4[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_44 = result_reg_r_4[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_45 = result_reg_r_4[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_46 = result_reg_r_4[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_47 = result_reg_r_4[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_48 = result_reg_r_4[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_49 = result_reg_r_4[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_50 = result_reg_r_4[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_51 = result_reg_r_4[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_52 = result_reg_r_4[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_53 = result_reg_r_4[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_54 = result_reg_r_4[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_55 = result_reg_r_4[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_56 = result_reg_r_4[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_57 = result_reg_r_4[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_58 = result_reg_r_4[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_59 = result_reg_r_4[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_60 = result_reg_r_4[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_61 = result_reg_r_4[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_62 = result_reg_r_4[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_63 = result_reg_r_4[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_64 = result_reg_r_4[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_65 = result_reg_r_4[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_66 = result_reg_r_4[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_67 = result_reg_r_4[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_68 = result_reg_r_4[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_69 = result_reg_r_4[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_70 = result_reg_r_4[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_71 = result_reg_r_4[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_72 = result_reg_r_4[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_73 = result_reg_r_4[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_74 = result_reg_r_4[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_75 = result_reg_r_4[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_76 = result_reg_r_4[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_77 = result_reg_r_4[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_78 = result_reg_r_4[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_79 = result_reg_r_4[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_80 = result_reg_r_4[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_81 = result_reg_r_4[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_82 = result_reg_r_4[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_83 = result_reg_r_4[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_84 = result_reg_r_4[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_85 = result_reg_r_4[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_86 = result_reg_r_4[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_87 = result_reg_r_4[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_88 = result_reg_r_4[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_89 = result_reg_r_4[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_90 = result_reg_r_4[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_91 = result_reg_r_4[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_92 = result_reg_r_4[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_93 = result_reg_r_4[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_94 = result_reg_r_4[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_96 = result_reg_r_4[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_97 = result_reg_r_4[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_98 = result_reg_r_4[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_99 = result_reg_r_4[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_100 = result_reg_r_4[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_101 = result_reg_r_4[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_102 = result_reg_r_4[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_103 = result_reg_r_4[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_104 = result_reg_r_4[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_9_105 = result_reg_r_4[105]; // @[BinaryDesigns2.scala 192:62]
  wire [200:0] _T_11256 = {b_aux_reg_r_4, 95'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [200:0] _GEN_1276 = {{95'd0}, a_aux_reg_r_4}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_9_95 = _GEN_1276 >= _T_11256; // @[BinaryDesigns2.scala 224:35]
  wire [6:0] result_reg_w_5_hi_hi_hi_lo = {wire_res_9_98,wire_res_9_97,wire_res_9_96,wire_res_9_95,wire_res_9_94,
    wire_res_9_93,wire_res_9_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_5_hi_hi_lo_lo = {wire_res_9_84,wire_res_9_83,wire_res_9_82,wire_res_9_81,wire_res_9_80,
    wire_res_9_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_5_hi_hi_lo = {wire_res_9_91,wire_res_9_90,wire_res_9_89,wire_res_9_88,wire_res_9_87,
    wire_res_9_86,wire_res_9_85,result_reg_w_5_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_5_hi_lo_hi_lo = {wire_res_9_71,wire_res_9_70,wire_res_9_69,wire_res_9_68,wire_res_9_67,
    wire_res_9_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_5_hi_lo_lo_lo = {wire_res_9_58,wire_res_9_57,wire_res_9_56,wire_res_9_55,wire_res_9_54,
    wire_res_9_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_5_hi_lo_lo = {wire_res_9_65,wire_res_9_64,wire_res_9_63,wire_res_9_62,wire_res_9_61,
    wire_res_9_60,wire_res_9_59,result_reg_w_5_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_5_hi_lo = {wire_res_9_78,wire_res_9_77,wire_res_9_76,wire_res_9_75,wire_res_9_74,
    wire_res_9_73,wire_res_9_72,result_reg_w_5_hi_lo_hi_lo,result_reg_w_5_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_5_hi = {wire_res_9_105,wire_res_9_104,wire_res_9_103,wire_res_9_102,wire_res_9_101,
    wire_res_9_100,wire_res_9_99,result_reg_w_5_hi_hi_hi_lo,result_reg_w_5_hi_hi_lo,result_reg_w_5_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_5_lo_hi_hi_lo = {wire_res_9_45,wire_res_9_44,wire_res_9_43,wire_res_9_42,wire_res_9_41,
    wire_res_9_40,wire_res_9_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_5_lo_hi_lo_lo = {wire_res_9_31,wire_res_9_30,wire_res_9_29,wire_res_9_28,wire_res_9_27,
    wire_res_9_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_5_lo_hi_lo = {wire_res_9_38,wire_res_9_37,wire_res_9_36,wire_res_9_35,wire_res_9_34,
    wire_res_9_33,wire_res_9_32,result_reg_w_5_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_5_lo_lo_hi_lo = {wire_res_9_18,wire_res_9_17,wire_res_9_16,wire_res_9_15,wire_res_9_14,
    wire_res_9_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_5_lo_lo_lo_lo = {wire_res_9_5,wire_res_9_4,wire_res_9_3,wire_res_9_2,wire_res_9_1,wire_res_9_0
    }; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_5_lo_lo_lo = {wire_res_9_12,wire_res_9_11,wire_res_9_10,wire_res_9_9,wire_res_9_8,
    wire_res_9_7,wire_res_9_6,result_reg_w_5_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_5_lo_lo = {wire_res_9_25,wire_res_9_24,wire_res_9_23,wire_res_9_22,wire_res_9_21,
    wire_res_9_20,wire_res_9_19,result_reg_w_5_lo_lo_hi_lo,result_reg_w_5_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_5_lo = {wire_res_9_52,wire_res_9_51,wire_res_9_50,wire_res_9_49,wire_res_9_48,wire_res_9_47,
    wire_res_9_46,result_reg_w_5_lo_hi_hi_lo,result_reg_w_5_lo_hi_lo,result_reg_w_5_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_5 = {result_reg_w_5_hi,result_reg_w_5_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_10_0 = result_reg_w_5[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_1 = result_reg_w_5[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_2 = result_reg_w_5[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_3 = result_reg_w_5[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_4 = result_reg_w_5[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_5 = result_reg_w_5[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_6 = result_reg_w_5[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_7 = result_reg_w_5[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_8 = result_reg_w_5[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_9 = result_reg_w_5[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_10 = result_reg_w_5[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_11 = result_reg_w_5[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_12 = result_reg_w_5[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_13 = result_reg_w_5[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_14 = result_reg_w_5[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_15 = result_reg_w_5[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_16 = result_reg_w_5[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_17 = result_reg_w_5[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_18 = result_reg_w_5[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_19 = result_reg_w_5[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_20 = result_reg_w_5[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_21 = result_reg_w_5[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_22 = result_reg_w_5[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_23 = result_reg_w_5[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_24 = result_reg_w_5[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_25 = result_reg_w_5[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_26 = result_reg_w_5[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_27 = result_reg_w_5[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_28 = result_reg_w_5[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_29 = result_reg_w_5[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_30 = result_reg_w_5[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_31 = result_reg_w_5[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_32 = result_reg_w_5[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_33 = result_reg_w_5[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_34 = result_reg_w_5[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_35 = result_reg_w_5[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_36 = result_reg_w_5[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_37 = result_reg_w_5[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_38 = result_reg_w_5[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_39 = result_reg_w_5[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_40 = result_reg_w_5[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_41 = result_reg_w_5[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_42 = result_reg_w_5[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_43 = result_reg_w_5[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_44 = result_reg_w_5[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_45 = result_reg_w_5[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_46 = result_reg_w_5[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_47 = result_reg_w_5[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_48 = result_reg_w_5[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_49 = result_reg_w_5[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_50 = result_reg_w_5[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_51 = result_reg_w_5[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_52 = result_reg_w_5[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_53 = result_reg_w_5[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_54 = result_reg_w_5[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_55 = result_reg_w_5[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_56 = result_reg_w_5[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_57 = result_reg_w_5[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_58 = result_reg_w_5[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_59 = result_reg_w_5[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_60 = result_reg_w_5[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_61 = result_reg_w_5[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_62 = result_reg_w_5[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_63 = result_reg_w_5[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_64 = result_reg_w_5[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_65 = result_reg_w_5[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_66 = result_reg_w_5[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_67 = result_reg_w_5[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_68 = result_reg_w_5[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_69 = result_reg_w_5[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_70 = result_reg_w_5[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_71 = result_reg_w_5[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_72 = result_reg_w_5[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_73 = result_reg_w_5[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_74 = result_reg_w_5[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_75 = result_reg_w_5[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_76 = result_reg_w_5[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_77 = result_reg_w_5[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_78 = result_reg_w_5[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_79 = result_reg_w_5[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_80 = result_reg_w_5[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_81 = result_reg_w_5[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_82 = result_reg_w_5[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_83 = result_reg_w_5[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_84 = result_reg_w_5[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_85 = result_reg_w_5[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_86 = result_reg_w_5[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_87 = result_reg_w_5[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_88 = result_reg_w_5[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_89 = result_reg_w_5[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_90 = result_reg_w_5[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_91 = result_reg_w_5[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_92 = result_reg_w_5[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_93 = result_reg_w_5[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_95 = result_reg_w_5[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_96 = result_reg_w_5[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_97 = result_reg_w_5[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_98 = result_reg_w_5[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_99 = result_reg_w_5[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_100 = result_reg_w_5[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_101 = result_reg_w_5[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_102 = result_reg_w_5[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_103 = result_reg_w_5[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_104 = result_reg_w_5[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_10_105 = result_reg_w_5[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_0 = result_reg_r_5[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_1 = result_reg_r_5[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_2 = result_reg_r_5[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_3 = result_reg_r_5[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_4 = result_reg_r_5[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_5 = result_reg_r_5[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_6 = result_reg_r_5[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_7 = result_reg_r_5[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_8 = result_reg_r_5[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_9 = result_reg_r_5[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_10 = result_reg_r_5[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_11 = result_reg_r_5[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_12 = result_reg_r_5[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_13 = result_reg_r_5[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_14 = result_reg_r_5[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_15 = result_reg_r_5[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_16 = result_reg_r_5[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_17 = result_reg_r_5[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_18 = result_reg_r_5[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_19 = result_reg_r_5[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_20 = result_reg_r_5[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_21 = result_reg_r_5[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_22 = result_reg_r_5[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_23 = result_reg_r_5[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_24 = result_reg_r_5[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_25 = result_reg_r_5[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_26 = result_reg_r_5[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_27 = result_reg_r_5[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_28 = result_reg_r_5[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_29 = result_reg_r_5[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_30 = result_reg_r_5[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_31 = result_reg_r_5[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_32 = result_reg_r_5[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_33 = result_reg_r_5[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_34 = result_reg_r_5[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_35 = result_reg_r_5[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_36 = result_reg_r_5[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_37 = result_reg_r_5[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_38 = result_reg_r_5[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_39 = result_reg_r_5[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_40 = result_reg_r_5[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_41 = result_reg_r_5[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_42 = result_reg_r_5[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_43 = result_reg_r_5[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_44 = result_reg_r_5[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_45 = result_reg_r_5[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_46 = result_reg_r_5[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_47 = result_reg_r_5[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_48 = result_reg_r_5[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_49 = result_reg_r_5[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_50 = result_reg_r_5[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_51 = result_reg_r_5[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_52 = result_reg_r_5[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_53 = result_reg_r_5[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_54 = result_reg_r_5[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_55 = result_reg_r_5[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_56 = result_reg_r_5[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_57 = result_reg_r_5[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_58 = result_reg_r_5[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_59 = result_reg_r_5[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_60 = result_reg_r_5[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_61 = result_reg_r_5[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_62 = result_reg_r_5[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_63 = result_reg_r_5[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_64 = result_reg_r_5[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_65 = result_reg_r_5[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_66 = result_reg_r_5[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_67 = result_reg_r_5[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_68 = result_reg_r_5[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_69 = result_reg_r_5[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_70 = result_reg_r_5[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_71 = result_reg_r_5[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_72 = result_reg_r_5[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_73 = result_reg_r_5[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_74 = result_reg_r_5[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_75 = result_reg_r_5[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_76 = result_reg_r_5[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_77 = result_reg_r_5[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_78 = result_reg_r_5[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_79 = result_reg_r_5[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_80 = result_reg_r_5[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_81 = result_reg_r_5[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_82 = result_reg_r_5[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_83 = result_reg_r_5[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_84 = result_reg_r_5[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_85 = result_reg_r_5[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_86 = result_reg_r_5[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_87 = result_reg_r_5[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_88 = result_reg_r_5[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_89 = result_reg_r_5[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_90 = result_reg_r_5[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_91 = result_reg_r_5[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_92 = result_reg_r_5[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_94 = result_reg_r_5[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_95 = result_reg_r_5[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_96 = result_reg_r_5[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_97 = result_reg_r_5[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_98 = result_reg_r_5[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_99 = result_reg_r_5[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_100 = result_reg_r_5[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_101 = result_reg_r_5[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_102 = result_reg_r_5[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_103 = result_reg_r_5[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_104 = result_reg_r_5[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_11_105 = result_reg_r_5[105]; // @[BinaryDesigns2.scala 192:62]
  wire [198:0] _T_11260 = {b_aux_reg_r_5, 93'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [198:0] _GEN_1277 = {{93'd0}, a_aux_reg_r_5}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_11_93 = _GEN_1277 >= _T_11260; // @[BinaryDesigns2.scala 224:35]
  wire [6:0] result_reg_w_6_hi_hi_hi_lo = {wire_res_11_98,wire_res_11_97,wire_res_11_96,wire_res_11_95,wire_res_11_94,
    wire_res_11_93,wire_res_11_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_6_hi_hi_lo_lo = {wire_res_11_84,wire_res_11_83,wire_res_11_82,wire_res_11_81,wire_res_11_80,
    wire_res_11_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_6_hi_hi_lo = {wire_res_11_91,wire_res_11_90,wire_res_11_89,wire_res_11_88,wire_res_11_87,
    wire_res_11_86,wire_res_11_85,result_reg_w_6_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_6_hi_lo_hi_lo = {wire_res_11_71,wire_res_11_70,wire_res_11_69,wire_res_11_68,wire_res_11_67,
    wire_res_11_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_6_hi_lo_lo_lo = {wire_res_11_58,wire_res_11_57,wire_res_11_56,wire_res_11_55,wire_res_11_54,
    wire_res_11_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_6_hi_lo_lo = {wire_res_11_65,wire_res_11_64,wire_res_11_63,wire_res_11_62,wire_res_11_61,
    wire_res_11_60,wire_res_11_59,result_reg_w_6_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_6_hi_lo = {wire_res_11_78,wire_res_11_77,wire_res_11_76,wire_res_11_75,wire_res_11_74,
    wire_res_11_73,wire_res_11_72,result_reg_w_6_hi_lo_hi_lo,result_reg_w_6_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_6_hi = {wire_res_11_105,wire_res_11_104,wire_res_11_103,wire_res_11_102,wire_res_11_101,
    wire_res_11_100,wire_res_11_99,result_reg_w_6_hi_hi_hi_lo,result_reg_w_6_hi_hi_lo,result_reg_w_6_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_6_lo_hi_hi_lo = {wire_res_11_45,wire_res_11_44,wire_res_11_43,wire_res_11_42,wire_res_11_41,
    wire_res_11_40,wire_res_11_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_6_lo_hi_lo_lo = {wire_res_11_31,wire_res_11_30,wire_res_11_29,wire_res_11_28,wire_res_11_27,
    wire_res_11_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_6_lo_hi_lo = {wire_res_11_38,wire_res_11_37,wire_res_11_36,wire_res_11_35,wire_res_11_34,
    wire_res_11_33,wire_res_11_32,result_reg_w_6_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_6_lo_lo_hi_lo = {wire_res_11_18,wire_res_11_17,wire_res_11_16,wire_res_11_15,wire_res_11_14,
    wire_res_11_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_6_lo_lo_lo_lo = {wire_res_11_5,wire_res_11_4,wire_res_11_3,wire_res_11_2,wire_res_11_1,
    wire_res_11_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_6_lo_lo_lo = {wire_res_11_12,wire_res_11_11,wire_res_11_10,wire_res_11_9,wire_res_11_8,
    wire_res_11_7,wire_res_11_6,result_reg_w_6_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_6_lo_lo = {wire_res_11_25,wire_res_11_24,wire_res_11_23,wire_res_11_22,wire_res_11_21,
    wire_res_11_20,wire_res_11_19,result_reg_w_6_lo_lo_hi_lo,result_reg_w_6_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_6_lo = {wire_res_11_52,wire_res_11_51,wire_res_11_50,wire_res_11_49,wire_res_11_48,
    wire_res_11_47,wire_res_11_46,result_reg_w_6_lo_hi_hi_lo,result_reg_w_6_lo_hi_lo,result_reg_w_6_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_6 = {result_reg_w_6_hi,result_reg_w_6_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_12_0 = result_reg_w_6[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_1 = result_reg_w_6[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_2 = result_reg_w_6[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_3 = result_reg_w_6[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_4 = result_reg_w_6[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_5 = result_reg_w_6[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_6 = result_reg_w_6[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_7 = result_reg_w_6[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_8 = result_reg_w_6[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_9 = result_reg_w_6[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_10 = result_reg_w_6[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_11 = result_reg_w_6[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_12 = result_reg_w_6[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_13 = result_reg_w_6[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_14 = result_reg_w_6[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_15 = result_reg_w_6[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_16 = result_reg_w_6[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_17 = result_reg_w_6[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_18 = result_reg_w_6[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_19 = result_reg_w_6[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_20 = result_reg_w_6[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_21 = result_reg_w_6[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_22 = result_reg_w_6[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_23 = result_reg_w_6[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_24 = result_reg_w_6[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_25 = result_reg_w_6[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_26 = result_reg_w_6[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_27 = result_reg_w_6[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_28 = result_reg_w_6[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_29 = result_reg_w_6[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_30 = result_reg_w_6[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_31 = result_reg_w_6[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_32 = result_reg_w_6[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_33 = result_reg_w_6[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_34 = result_reg_w_6[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_35 = result_reg_w_6[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_36 = result_reg_w_6[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_37 = result_reg_w_6[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_38 = result_reg_w_6[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_39 = result_reg_w_6[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_40 = result_reg_w_6[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_41 = result_reg_w_6[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_42 = result_reg_w_6[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_43 = result_reg_w_6[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_44 = result_reg_w_6[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_45 = result_reg_w_6[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_46 = result_reg_w_6[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_47 = result_reg_w_6[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_48 = result_reg_w_6[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_49 = result_reg_w_6[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_50 = result_reg_w_6[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_51 = result_reg_w_6[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_52 = result_reg_w_6[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_53 = result_reg_w_6[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_54 = result_reg_w_6[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_55 = result_reg_w_6[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_56 = result_reg_w_6[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_57 = result_reg_w_6[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_58 = result_reg_w_6[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_59 = result_reg_w_6[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_60 = result_reg_w_6[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_61 = result_reg_w_6[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_62 = result_reg_w_6[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_63 = result_reg_w_6[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_64 = result_reg_w_6[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_65 = result_reg_w_6[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_66 = result_reg_w_6[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_67 = result_reg_w_6[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_68 = result_reg_w_6[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_69 = result_reg_w_6[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_70 = result_reg_w_6[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_71 = result_reg_w_6[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_72 = result_reg_w_6[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_73 = result_reg_w_6[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_74 = result_reg_w_6[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_75 = result_reg_w_6[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_76 = result_reg_w_6[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_77 = result_reg_w_6[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_78 = result_reg_w_6[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_79 = result_reg_w_6[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_80 = result_reg_w_6[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_81 = result_reg_w_6[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_82 = result_reg_w_6[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_83 = result_reg_w_6[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_84 = result_reg_w_6[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_85 = result_reg_w_6[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_86 = result_reg_w_6[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_87 = result_reg_w_6[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_88 = result_reg_w_6[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_89 = result_reg_w_6[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_90 = result_reg_w_6[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_91 = result_reg_w_6[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_93 = result_reg_w_6[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_94 = result_reg_w_6[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_95 = result_reg_w_6[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_96 = result_reg_w_6[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_97 = result_reg_w_6[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_98 = result_reg_w_6[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_99 = result_reg_w_6[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_100 = result_reg_w_6[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_101 = result_reg_w_6[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_102 = result_reg_w_6[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_103 = result_reg_w_6[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_104 = result_reg_w_6[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_12_105 = result_reg_w_6[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_0 = result_reg_r_6[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_1 = result_reg_r_6[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_2 = result_reg_r_6[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_3 = result_reg_r_6[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_4 = result_reg_r_6[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_5 = result_reg_r_6[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_6 = result_reg_r_6[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_7 = result_reg_r_6[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_8 = result_reg_r_6[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_9 = result_reg_r_6[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_10 = result_reg_r_6[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_11 = result_reg_r_6[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_12 = result_reg_r_6[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_13 = result_reg_r_6[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_14 = result_reg_r_6[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_15 = result_reg_r_6[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_16 = result_reg_r_6[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_17 = result_reg_r_6[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_18 = result_reg_r_6[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_19 = result_reg_r_6[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_20 = result_reg_r_6[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_21 = result_reg_r_6[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_22 = result_reg_r_6[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_23 = result_reg_r_6[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_24 = result_reg_r_6[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_25 = result_reg_r_6[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_26 = result_reg_r_6[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_27 = result_reg_r_6[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_28 = result_reg_r_6[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_29 = result_reg_r_6[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_30 = result_reg_r_6[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_31 = result_reg_r_6[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_32 = result_reg_r_6[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_33 = result_reg_r_6[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_34 = result_reg_r_6[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_35 = result_reg_r_6[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_36 = result_reg_r_6[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_37 = result_reg_r_6[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_38 = result_reg_r_6[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_39 = result_reg_r_6[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_40 = result_reg_r_6[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_41 = result_reg_r_6[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_42 = result_reg_r_6[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_43 = result_reg_r_6[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_44 = result_reg_r_6[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_45 = result_reg_r_6[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_46 = result_reg_r_6[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_47 = result_reg_r_6[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_48 = result_reg_r_6[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_49 = result_reg_r_6[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_50 = result_reg_r_6[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_51 = result_reg_r_6[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_52 = result_reg_r_6[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_53 = result_reg_r_6[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_54 = result_reg_r_6[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_55 = result_reg_r_6[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_56 = result_reg_r_6[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_57 = result_reg_r_6[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_58 = result_reg_r_6[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_59 = result_reg_r_6[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_60 = result_reg_r_6[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_61 = result_reg_r_6[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_62 = result_reg_r_6[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_63 = result_reg_r_6[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_64 = result_reg_r_6[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_65 = result_reg_r_6[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_66 = result_reg_r_6[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_67 = result_reg_r_6[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_68 = result_reg_r_6[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_69 = result_reg_r_6[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_70 = result_reg_r_6[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_71 = result_reg_r_6[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_72 = result_reg_r_6[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_73 = result_reg_r_6[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_74 = result_reg_r_6[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_75 = result_reg_r_6[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_76 = result_reg_r_6[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_77 = result_reg_r_6[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_78 = result_reg_r_6[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_79 = result_reg_r_6[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_80 = result_reg_r_6[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_81 = result_reg_r_6[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_82 = result_reg_r_6[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_83 = result_reg_r_6[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_84 = result_reg_r_6[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_85 = result_reg_r_6[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_86 = result_reg_r_6[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_87 = result_reg_r_6[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_88 = result_reg_r_6[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_89 = result_reg_r_6[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_90 = result_reg_r_6[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_92 = result_reg_r_6[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_93 = result_reg_r_6[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_94 = result_reg_r_6[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_95 = result_reg_r_6[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_96 = result_reg_r_6[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_97 = result_reg_r_6[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_98 = result_reg_r_6[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_99 = result_reg_r_6[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_100 = result_reg_r_6[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_101 = result_reg_r_6[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_102 = result_reg_r_6[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_103 = result_reg_r_6[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_104 = result_reg_r_6[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_13_105 = result_reg_r_6[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_7_hi_hi_hi_lo = {wire_res_13_98,wire_res_13_97,wire_res_13_96,wire_res_13_95,wire_res_13_94,
    wire_res_13_93,wire_res_13_92}; // @[BinaryDesigns2.scala 231:46]
  wire [196:0] _T_11264 = {b_aux_reg_r_6, 91'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [196:0] _GEN_1278 = {{91'd0}, a_aux_reg_r_6}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_13_91 = _GEN_1278 >= _T_11264; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_7_hi_hi_lo_lo = {wire_res_13_84,wire_res_13_83,wire_res_13_82,wire_res_13_81,wire_res_13_80,
    wire_res_13_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_7_hi_hi_lo = {wire_res_13_91,wire_res_13_90,wire_res_13_89,wire_res_13_88,wire_res_13_87,
    wire_res_13_86,wire_res_13_85,result_reg_w_7_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_7_hi_lo_hi_lo = {wire_res_13_71,wire_res_13_70,wire_res_13_69,wire_res_13_68,wire_res_13_67,
    wire_res_13_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_7_hi_lo_lo_lo = {wire_res_13_58,wire_res_13_57,wire_res_13_56,wire_res_13_55,wire_res_13_54,
    wire_res_13_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_7_hi_lo_lo = {wire_res_13_65,wire_res_13_64,wire_res_13_63,wire_res_13_62,wire_res_13_61,
    wire_res_13_60,wire_res_13_59,result_reg_w_7_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_7_hi_lo = {wire_res_13_78,wire_res_13_77,wire_res_13_76,wire_res_13_75,wire_res_13_74,
    wire_res_13_73,wire_res_13_72,result_reg_w_7_hi_lo_hi_lo,result_reg_w_7_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_7_hi = {wire_res_13_105,wire_res_13_104,wire_res_13_103,wire_res_13_102,wire_res_13_101,
    wire_res_13_100,wire_res_13_99,result_reg_w_7_hi_hi_hi_lo,result_reg_w_7_hi_hi_lo,result_reg_w_7_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_7_lo_hi_hi_lo = {wire_res_13_45,wire_res_13_44,wire_res_13_43,wire_res_13_42,wire_res_13_41,
    wire_res_13_40,wire_res_13_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_7_lo_hi_lo_lo = {wire_res_13_31,wire_res_13_30,wire_res_13_29,wire_res_13_28,wire_res_13_27,
    wire_res_13_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_7_lo_hi_lo = {wire_res_13_38,wire_res_13_37,wire_res_13_36,wire_res_13_35,wire_res_13_34,
    wire_res_13_33,wire_res_13_32,result_reg_w_7_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_7_lo_lo_hi_lo = {wire_res_13_18,wire_res_13_17,wire_res_13_16,wire_res_13_15,wire_res_13_14,
    wire_res_13_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_7_lo_lo_lo_lo = {wire_res_13_5,wire_res_13_4,wire_res_13_3,wire_res_13_2,wire_res_13_1,
    wire_res_13_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_7_lo_lo_lo = {wire_res_13_12,wire_res_13_11,wire_res_13_10,wire_res_13_9,wire_res_13_8,
    wire_res_13_7,wire_res_13_6,result_reg_w_7_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_7_lo_lo = {wire_res_13_25,wire_res_13_24,wire_res_13_23,wire_res_13_22,wire_res_13_21,
    wire_res_13_20,wire_res_13_19,result_reg_w_7_lo_lo_hi_lo,result_reg_w_7_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_7_lo = {wire_res_13_52,wire_res_13_51,wire_res_13_50,wire_res_13_49,wire_res_13_48,
    wire_res_13_47,wire_res_13_46,result_reg_w_7_lo_hi_hi_lo,result_reg_w_7_lo_hi_lo,result_reg_w_7_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_7 = {result_reg_w_7_hi,result_reg_w_7_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_14_0 = result_reg_w_7[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_1 = result_reg_w_7[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_2 = result_reg_w_7[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_3 = result_reg_w_7[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_4 = result_reg_w_7[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_5 = result_reg_w_7[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_6 = result_reg_w_7[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_7 = result_reg_w_7[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_8 = result_reg_w_7[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_9 = result_reg_w_7[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_10 = result_reg_w_7[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_11 = result_reg_w_7[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_12 = result_reg_w_7[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_13 = result_reg_w_7[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_14 = result_reg_w_7[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_15 = result_reg_w_7[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_16 = result_reg_w_7[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_17 = result_reg_w_7[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_18 = result_reg_w_7[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_19 = result_reg_w_7[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_20 = result_reg_w_7[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_21 = result_reg_w_7[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_22 = result_reg_w_7[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_23 = result_reg_w_7[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_24 = result_reg_w_7[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_25 = result_reg_w_7[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_26 = result_reg_w_7[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_27 = result_reg_w_7[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_28 = result_reg_w_7[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_29 = result_reg_w_7[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_30 = result_reg_w_7[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_31 = result_reg_w_7[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_32 = result_reg_w_7[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_33 = result_reg_w_7[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_34 = result_reg_w_7[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_35 = result_reg_w_7[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_36 = result_reg_w_7[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_37 = result_reg_w_7[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_38 = result_reg_w_7[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_39 = result_reg_w_7[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_40 = result_reg_w_7[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_41 = result_reg_w_7[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_42 = result_reg_w_7[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_43 = result_reg_w_7[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_44 = result_reg_w_7[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_45 = result_reg_w_7[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_46 = result_reg_w_7[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_47 = result_reg_w_7[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_48 = result_reg_w_7[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_49 = result_reg_w_7[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_50 = result_reg_w_7[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_51 = result_reg_w_7[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_52 = result_reg_w_7[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_53 = result_reg_w_7[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_54 = result_reg_w_7[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_55 = result_reg_w_7[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_56 = result_reg_w_7[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_57 = result_reg_w_7[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_58 = result_reg_w_7[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_59 = result_reg_w_7[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_60 = result_reg_w_7[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_61 = result_reg_w_7[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_62 = result_reg_w_7[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_63 = result_reg_w_7[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_64 = result_reg_w_7[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_65 = result_reg_w_7[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_66 = result_reg_w_7[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_67 = result_reg_w_7[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_68 = result_reg_w_7[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_69 = result_reg_w_7[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_70 = result_reg_w_7[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_71 = result_reg_w_7[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_72 = result_reg_w_7[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_73 = result_reg_w_7[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_74 = result_reg_w_7[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_75 = result_reg_w_7[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_76 = result_reg_w_7[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_77 = result_reg_w_7[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_78 = result_reg_w_7[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_79 = result_reg_w_7[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_80 = result_reg_w_7[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_81 = result_reg_w_7[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_82 = result_reg_w_7[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_83 = result_reg_w_7[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_84 = result_reg_w_7[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_85 = result_reg_w_7[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_86 = result_reg_w_7[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_87 = result_reg_w_7[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_88 = result_reg_w_7[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_89 = result_reg_w_7[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_91 = result_reg_w_7[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_92 = result_reg_w_7[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_93 = result_reg_w_7[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_94 = result_reg_w_7[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_95 = result_reg_w_7[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_96 = result_reg_w_7[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_97 = result_reg_w_7[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_98 = result_reg_w_7[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_99 = result_reg_w_7[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_100 = result_reg_w_7[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_101 = result_reg_w_7[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_102 = result_reg_w_7[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_103 = result_reg_w_7[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_104 = result_reg_w_7[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_14_105 = result_reg_w_7[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_0 = result_reg_r_7[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_1 = result_reg_r_7[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_2 = result_reg_r_7[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_3 = result_reg_r_7[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_4 = result_reg_r_7[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_5 = result_reg_r_7[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_6 = result_reg_r_7[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_7 = result_reg_r_7[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_8 = result_reg_r_7[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_9 = result_reg_r_7[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_10 = result_reg_r_7[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_11 = result_reg_r_7[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_12 = result_reg_r_7[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_13 = result_reg_r_7[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_14 = result_reg_r_7[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_15 = result_reg_r_7[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_16 = result_reg_r_7[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_17 = result_reg_r_7[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_18 = result_reg_r_7[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_19 = result_reg_r_7[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_20 = result_reg_r_7[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_21 = result_reg_r_7[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_22 = result_reg_r_7[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_23 = result_reg_r_7[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_24 = result_reg_r_7[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_25 = result_reg_r_7[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_26 = result_reg_r_7[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_27 = result_reg_r_7[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_28 = result_reg_r_7[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_29 = result_reg_r_7[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_30 = result_reg_r_7[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_31 = result_reg_r_7[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_32 = result_reg_r_7[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_33 = result_reg_r_7[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_34 = result_reg_r_7[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_35 = result_reg_r_7[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_36 = result_reg_r_7[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_37 = result_reg_r_7[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_38 = result_reg_r_7[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_39 = result_reg_r_7[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_40 = result_reg_r_7[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_41 = result_reg_r_7[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_42 = result_reg_r_7[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_43 = result_reg_r_7[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_44 = result_reg_r_7[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_45 = result_reg_r_7[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_46 = result_reg_r_7[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_47 = result_reg_r_7[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_48 = result_reg_r_7[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_49 = result_reg_r_7[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_50 = result_reg_r_7[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_51 = result_reg_r_7[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_52 = result_reg_r_7[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_53 = result_reg_r_7[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_54 = result_reg_r_7[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_55 = result_reg_r_7[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_56 = result_reg_r_7[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_57 = result_reg_r_7[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_58 = result_reg_r_7[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_59 = result_reg_r_7[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_60 = result_reg_r_7[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_61 = result_reg_r_7[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_62 = result_reg_r_7[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_63 = result_reg_r_7[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_64 = result_reg_r_7[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_65 = result_reg_r_7[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_66 = result_reg_r_7[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_67 = result_reg_r_7[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_68 = result_reg_r_7[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_69 = result_reg_r_7[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_70 = result_reg_r_7[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_71 = result_reg_r_7[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_72 = result_reg_r_7[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_73 = result_reg_r_7[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_74 = result_reg_r_7[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_75 = result_reg_r_7[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_76 = result_reg_r_7[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_77 = result_reg_r_7[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_78 = result_reg_r_7[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_79 = result_reg_r_7[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_80 = result_reg_r_7[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_81 = result_reg_r_7[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_82 = result_reg_r_7[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_83 = result_reg_r_7[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_84 = result_reg_r_7[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_85 = result_reg_r_7[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_86 = result_reg_r_7[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_87 = result_reg_r_7[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_88 = result_reg_r_7[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_90 = result_reg_r_7[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_91 = result_reg_r_7[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_92 = result_reg_r_7[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_93 = result_reg_r_7[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_94 = result_reg_r_7[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_95 = result_reg_r_7[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_96 = result_reg_r_7[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_97 = result_reg_r_7[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_98 = result_reg_r_7[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_99 = result_reg_r_7[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_100 = result_reg_r_7[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_101 = result_reg_r_7[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_102 = result_reg_r_7[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_103 = result_reg_r_7[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_104 = result_reg_r_7[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_15_105 = result_reg_r_7[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_8_hi_hi_hi_lo = {wire_res_15_98,wire_res_15_97,wire_res_15_96,wire_res_15_95,wire_res_15_94,
    wire_res_15_93,wire_res_15_92}; // @[BinaryDesigns2.scala 231:46]
  wire [194:0] _T_11268 = {b_aux_reg_r_7, 89'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [194:0] _GEN_1279 = {{89'd0}, a_aux_reg_r_7}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_15_89 = _GEN_1279 >= _T_11268; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_8_hi_hi_lo_lo = {wire_res_15_84,wire_res_15_83,wire_res_15_82,wire_res_15_81,wire_res_15_80,
    wire_res_15_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_8_hi_hi_lo = {wire_res_15_91,wire_res_15_90,wire_res_15_89,wire_res_15_88,wire_res_15_87,
    wire_res_15_86,wire_res_15_85,result_reg_w_8_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_8_hi_lo_hi_lo = {wire_res_15_71,wire_res_15_70,wire_res_15_69,wire_res_15_68,wire_res_15_67,
    wire_res_15_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_8_hi_lo_lo_lo = {wire_res_15_58,wire_res_15_57,wire_res_15_56,wire_res_15_55,wire_res_15_54,
    wire_res_15_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_8_hi_lo_lo = {wire_res_15_65,wire_res_15_64,wire_res_15_63,wire_res_15_62,wire_res_15_61,
    wire_res_15_60,wire_res_15_59,result_reg_w_8_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_8_hi_lo = {wire_res_15_78,wire_res_15_77,wire_res_15_76,wire_res_15_75,wire_res_15_74,
    wire_res_15_73,wire_res_15_72,result_reg_w_8_hi_lo_hi_lo,result_reg_w_8_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_8_hi = {wire_res_15_105,wire_res_15_104,wire_res_15_103,wire_res_15_102,wire_res_15_101,
    wire_res_15_100,wire_res_15_99,result_reg_w_8_hi_hi_hi_lo,result_reg_w_8_hi_hi_lo,result_reg_w_8_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_8_lo_hi_hi_lo = {wire_res_15_45,wire_res_15_44,wire_res_15_43,wire_res_15_42,wire_res_15_41,
    wire_res_15_40,wire_res_15_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_8_lo_hi_lo_lo = {wire_res_15_31,wire_res_15_30,wire_res_15_29,wire_res_15_28,wire_res_15_27,
    wire_res_15_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_8_lo_hi_lo = {wire_res_15_38,wire_res_15_37,wire_res_15_36,wire_res_15_35,wire_res_15_34,
    wire_res_15_33,wire_res_15_32,result_reg_w_8_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_8_lo_lo_hi_lo = {wire_res_15_18,wire_res_15_17,wire_res_15_16,wire_res_15_15,wire_res_15_14,
    wire_res_15_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_8_lo_lo_lo_lo = {wire_res_15_5,wire_res_15_4,wire_res_15_3,wire_res_15_2,wire_res_15_1,
    wire_res_15_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_8_lo_lo_lo = {wire_res_15_12,wire_res_15_11,wire_res_15_10,wire_res_15_9,wire_res_15_8,
    wire_res_15_7,wire_res_15_6,result_reg_w_8_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_8_lo_lo = {wire_res_15_25,wire_res_15_24,wire_res_15_23,wire_res_15_22,wire_res_15_21,
    wire_res_15_20,wire_res_15_19,result_reg_w_8_lo_lo_hi_lo,result_reg_w_8_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_8_lo = {wire_res_15_52,wire_res_15_51,wire_res_15_50,wire_res_15_49,wire_res_15_48,
    wire_res_15_47,wire_res_15_46,result_reg_w_8_lo_hi_hi_lo,result_reg_w_8_lo_hi_lo,result_reg_w_8_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_8 = {result_reg_w_8_hi,result_reg_w_8_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_16_0 = result_reg_w_8[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_1 = result_reg_w_8[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_2 = result_reg_w_8[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_3 = result_reg_w_8[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_4 = result_reg_w_8[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_5 = result_reg_w_8[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_6 = result_reg_w_8[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_7 = result_reg_w_8[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_8 = result_reg_w_8[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_9 = result_reg_w_8[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_10 = result_reg_w_8[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_11 = result_reg_w_8[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_12 = result_reg_w_8[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_13 = result_reg_w_8[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_14 = result_reg_w_8[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_15 = result_reg_w_8[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_16 = result_reg_w_8[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_17 = result_reg_w_8[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_18 = result_reg_w_8[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_19 = result_reg_w_8[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_20 = result_reg_w_8[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_21 = result_reg_w_8[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_22 = result_reg_w_8[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_23 = result_reg_w_8[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_24 = result_reg_w_8[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_25 = result_reg_w_8[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_26 = result_reg_w_8[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_27 = result_reg_w_8[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_28 = result_reg_w_8[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_29 = result_reg_w_8[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_30 = result_reg_w_8[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_31 = result_reg_w_8[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_32 = result_reg_w_8[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_33 = result_reg_w_8[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_34 = result_reg_w_8[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_35 = result_reg_w_8[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_36 = result_reg_w_8[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_37 = result_reg_w_8[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_38 = result_reg_w_8[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_39 = result_reg_w_8[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_40 = result_reg_w_8[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_41 = result_reg_w_8[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_42 = result_reg_w_8[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_43 = result_reg_w_8[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_44 = result_reg_w_8[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_45 = result_reg_w_8[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_46 = result_reg_w_8[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_47 = result_reg_w_8[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_48 = result_reg_w_8[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_49 = result_reg_w_8[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_50 = result_reg_w_8[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_51 = result_reg_w_8[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_52 = result_reg_w_8[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_53 = result_reg_w_8[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_54 = result_reg_w_8[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_55 = result_reg_w_8[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_56 = result_reg_w_8[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_57 = result_reg_w_8[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_58 = result_reg_w_8[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_59 = result_reg_w_8[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_60 = result_reg_w_8[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_61 = result_reg_w_8[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_62 = result_reg_w_8[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_63 = result_reg_w_8[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_64 = result_reg_w_8[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_65 = result_reg_w_8[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_66 = result_reg_w_8[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_67 = result_reg_w_8[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_68 = result_reg_w_8[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_69 = result_reg_w_8[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_70 = result_reg_w_8[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_71 = result_reg_w_8[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_72 = result_reg_w_8[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_73 = result_reg_w_8[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_74 = result_reg_w_8[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_75 = result_reg_w_8[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_76 = result_reg_w_8[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_77 = result_reg_w_8[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_78 = result_reg_w_8[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_79 = result_reg_w_8[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_80 = result_reg_w_8[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_81 = result_reg_w_8[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_82 = result_reg_w_8[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_83 = result_reg_w_8[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_84 = result_reg_w_8[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_85 = result_reg_w_8[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_86 = result_reg_w_8[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_87 = result_reg_w_8[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_89 = result_reg_w_8[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_90 = result_reg_w_8[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_91 = result_reg_w_8[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_92 = result_reg_w_8[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_93 = result_reg_w_8[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_94 = result_reg_w_8[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_95 = result_reg_w_8[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_96 = result_reg_w_8[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_97 = result_reg_w_8[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_98 = result_reg_w_8[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_99 = result_reg_w_8[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_100 = result_reg_w_8[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_101 = result_reg_w_8[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_102 = result_reg_w_8[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_103 = result_reg_w_8[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_104 = result_reg_w_8[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_16_105 = result_reg_w_8[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_0 = result_reg_r_8[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_1 = result_reg_r_8[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_2 = result_reg_r_8[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_3 = result_reg_r_8[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_4 = result_reg_r_8[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_5 = result_reg_r_8[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_6 = result_reg_r_8[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_7 = result_reg_r_8[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_8 = result_reg_r_8[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_9 = result_reg_r_8[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_10 = result_reg_r_8[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_11 = result_reg_r_8[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_12 = result_reg_r_8[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_13 = result_reg_r_8[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_14 = result_reg_r_8[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_15 = result_reg_r_8[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_16 = result_reg_r_8[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_17 = result_reg_r_8[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_18 = result_reg_r_8[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_19 = result_reg_r_8[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_20 = result_reg_r_8[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_21 = result_reg_r_8[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_22 = result_reg_r_8[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_23 = result_reg_r_8[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_24 = result_reg_r_8[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_25 = result_reg_r_8[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_26 = result_reg_r_8[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_27 = result_reg_r_8[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_28 = result_reg_r_8[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_29 = result_reg_r_8[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_30 = result_reg_r_8[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_31 = result_reg_r_8[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_32 = result_reg_r_8[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_33 = result_reg_r_8[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_34 = result_reg_r_8[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_35 = result_reg_r_8[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_36 = result_reg_r_8[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_37 = result_reg_r_8[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_38 = result_reg_r_8[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_39 = result_reg_r_8[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_40 = result_reg_r_8[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_41 = result_reg_r_8[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_42 = result_reg_r_8[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_43 = result_reg_r_8[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_44 = result_reg_r_8[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_45 = result_reg_r_8[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_46 = result_reg_r_8[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_47 = result_reg_r_8[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_48 = result_reg_r_8[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_49 = result_reg_r_8[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_50 = result_reg_r_8[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_51 = result_reg_r_8[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_52 = result_reg_r_8[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_53 = result_reg_r_8[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_54 = result_reg_r_8[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_55 = result_reg_r_8[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_56 = result_reg_r_8[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_57 = result_reg_r_8[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_58 = result_reg_r_8[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_59 = result_reg_r_8[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_60 = result_reg_r_8[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_61 = result_reg_r_8[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_62 = result_reg_r_8[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_63 = result_reg_r_8[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_64 = result_reg_r_8[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_65 = result_reg_r_8[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_66 = result_reg_r_8[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_67 = result_reg_r_8[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_68 = result_reg_r_8[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_69 = result_reg_r_8[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_70 = result_reg_r_8[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_71 = result_reg_r_8[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_72 = result_reg_r_8[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_73 = result_reg_r_8[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_74 = result_reg_r_8[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_75 = result_reg_r_8[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_76 = result_reg_r_8[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_77 = result_reg_r_8[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_78 = result_reg_r_8[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_79 = result_reg_r_8[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_80 = result_reg_r_8[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_81 = result_reg_r_8[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_82 = result_reg_r_8[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_83 = result_reg_r_8[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_84 = result_reg_r_8[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_85 = result_reg_r_8[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_86 = result_reg_r_8[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_88 = result_reg_r_8[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_89 = result_reg_r_8[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_90 = result_reg_r_8[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_91 = result_reg_r_8[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_92 = result_reg_r_8[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_93 = result_reg_r_8[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_94 = result_reg_r_8[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_95 = result_reg_r_8[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_96 = result_reg_r_8[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_97 = result_reg_r_8[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_98 = result_reg_r_8[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_99 = result_reg_r_8[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_100 = result_reg_r_8[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_101 = result_reg_r_8[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_102 = result_reg_r_8[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_103 = result_reg_r_8[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_104 = result_reg_r_8[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_17_105 = result_reg_r_8[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_9_hi_hi_hi_lo = {wire_res_17_98,wire_res_17_97,wire_res_17_96,wire_res_17_95,wire_res_17_94,
    wire_res_17_93,wire_res_17_92}; // @[BinaryDesigns2.scala 231:46]
  wire [192:0] _T_11272 = {b_aux_reg_r_8, 87'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [192:0] _GEN_1280 = {{87'd0}, a_aux_reg_r_8}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_17_87 = _GEN_1280 >= _T_11272; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_9_hi_hi_lo_lo = {wire_res_17_84,wire_res_17_83,wire_res_17_82,wire_res_17_81,wire_res_17_80,
    wire_res_17_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_9_hi_hi_lo = {wire_res_17_91,wire_res_17_90,wire_res_17_89,wire_res_17_88,wire_res_17_87,
    wire_res_17_86,wire_res_17_85,result_reg_w_9_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_9_hi_lo_hi_lo = {wire_res_17_71,wire_res_17_70,wire_res_17_69,wire_res_17_68,wire_res_17_67,
    wire_res_17_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_9_hi_lo_lo_lo = {wire_res_17_58,wire_res_17_57,wire_res_17_56,wire_res_17_55,wire_res_17_54,
    wire_res_17_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_9_hi_lo_lo = {wire_res_17_65,wire_res_17_64,wire_res_17_63,wire_res_17_62,wire_res_17_61,
    wire_res_17_60,wire_res_17_59,result_reg_w_9_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_9_hi_lo = {wire_res_17_78,wire_res_17_77,wire_res_17_76,wire_res_17_75,wire_res_17_74,
    wire_res_17_73,wire_res_17_72,result_reg_w_9_hi_lo_hi_lo,result_reg_w_9_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_9_hi = {wire_res_17_105,wire_res_17_104,wire_res_17_103,wire_res_17_102,wire_res_17_101,
    wire_res_17_100,wire_res_17_99,result_reg_w_9_hi_hi_hi_lo,result_reg_w_9_hi_hi_lo,result_reg_w_9_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_9_lo_hi_hi_lo = {wire_res_17_45,wire_res_17_44,wire_res_17_43,wire_res_17_42,wire_res_17_41,
    wire_res_17_40,wire_res_17_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_9_lo_hi_lo_lo = {wire_res_17_31,wire_res_17_30,wire_res_17_29,wire_res_17_28,wire_res_17_27,
    wire_res_17_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_9_lo_hi_lo = {wire_res_17_38,wire_res_17_37,wire_res_17_36,wire_res_17_35,wire_res_17_34,
    wire_res_17_33,wire_res_17_32,result_reg_w_9_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_9_lo_lo_hi_lo = {wire_res_17_18,wire_res_17_17,wire_res_17_16,wire_res_17_15,wire_res_17_14,
    wire_res_17_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_9_lo_lo_lo_lo = {wire_res_17_5,wire_res_17_4,wire_res_17_3,wire_res_17_2,wire_res_17_1,
    wire_res_17_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_9_lo_lo_lo = {wire_res_17_12,wire_res_17_11,wire_res_17_10,wire_res_17_9,wire_res_17_8,
    wire_res_17_7,wire_res_17_6,result_reg_w_9_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_9_lo_lo = {wire_res_17_25,wire_res_17_24,wire_res_17_23,wire_res_17_22,wire_res_17_21,
    wire_res_17_20,wire_res_17_19,result_reg_w_9_lo_lo_hi_lo,result_reg_w_9_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_9_lo = {wire_res_17_52,wire_res_17_51,wire_res_17_50,wire_res_17_49,wire_res_17_48,
    wire_res_17_47,wire_res_17_46,result_reg_w_9_lo_hi_hi_lo,result_reg_w_9_lo_hi_lo,result_reg_w_9_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_9 = {result_reg_w_9_hi,result_reg_w_9_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_18_0 = result_reg_w_9[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_1 = result_reg_w_9[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_2 = result_reg_w_9[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_3 = result_reg_w_9[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_4 = result_reg_w_9[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_5 = result_reg_w_9[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_6 = result_reg_w_9[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_7 = result_reg_w_9[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_8 = result_reg_w_9[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_9 = result_reg_w_9[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_10 = result_reg_w_9[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_11 = result_reg_w_9[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_12 = result_reg_w_9[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_13 = result_reg_w_9[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_14 = result_reg_w_9[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_15 = result_reg_w_9[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_16 = result_reg_w_9[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_17 = result_reg_w_9[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_18 = result_reg_w_9[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_19 = result_reg_w_9[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_20 = result_reg_w_9[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_21 = result_reg_w_9[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_22 = result_reg_w_9[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_23 = result_reg_w_9[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_24 = result_reg_w_9[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_25 = result_reg_w_9[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_26 = result_reg_w_9[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_27 = result_reg_w_9[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_28 = result_reg_w_9[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_29 = result_reg_w_9[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_30 = result_reg_w_9[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_31 = result_reg_w_9[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_32 = result_reg_w_9[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_33 = result_reg_w_9[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_34 = result_reg_w_9[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_35 = result_reg_w_9[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_36 = result_reg_w_9[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_37 = result_reg_w_9[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_38 = result_reg_w_9[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_39 = result_reg_w_9[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_40 = result_reg_w_9[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_41 = result_reg_w_9[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_42 = result_reg_w_9[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_43 = result_reg_w_9[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_44 = result_reg_w_9[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_45 = result_reg_w_9[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_46 = result_reg_w_9[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_47 = result_reg_w_9[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_48 = result_reg_w_9[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_49 = result_reg_w_9[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_50 = result_reg_w_9[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_51 = result_reg_w_9[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_52 = result_reg_w_9[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_53 = result_reg_w_9[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_54 = result_reg_w_9[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_55 = result_reg_w_9[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_56 = result_reg_w_9[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_57 = result_reg_w_9[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_58 = result_reg_w_9[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_59 = result_reg_w_9[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_60 = result_reg_w_9[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_61 = result_reg_w_9[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_62 = result_reg_w_9[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_63 = result_reg_w_9[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_64 = result_reg_w_9[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_65 = result_reg_w_9[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_66 = result_reg_w_9[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_67 = result_reg_w_9[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_68 = result_reg_w_9[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_69 = result_reg_w_9[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_70 = result_reg_w_9[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_71 = result_reg_w_9[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_72 = result_reg_w_9[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_73 = result_reg_w_9[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_74 = result_reg_w_9[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_75 = result_reg_w_9[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_76 = result_reg_w_9[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_77 = result_reg_w_9[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_78 = result_reg_w_9[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_79 = result_reg_w_9[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_80 = result_reg_w_9[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_81 = result_reg_w_9[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_82 = result_reg_w_9[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_83 = result_reg_w_9[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_84 = result_reg_w_9[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_85 = result_reg_w_9[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_87 = result_reg_w_9[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_88 = result_reg_w_9[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_89 = result_reg_w_9[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_90 = result_reg_w_9[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_91 = result_reg_w_9[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_92 = result_reg_w_9[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_93 = result_reg_w_9[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_94 = result_reg_w_9[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_95 = result_reg_w_9[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_96 = result_reg_w_9[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_97 = result_reg_w_9[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_98 = result_reg_w_9[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_99 = result_reg_w_9[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_100 = result_reg_w_9[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_101 = result_reg_w_9[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_102 = result_reg_w_9[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_103 = result_reg_w_9[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_104 = result_reg_w_9[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_18_105 = result_reg_w_9[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_0 = result_reg_r_9[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_1 = result_reg_r_9[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_2 = result_reg_r_9[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_3 = result_reg_r_9[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_4 = result_reg_r_9[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_5 = result_reg_r_9[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_6 = result_reg_r_9[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_7 = result_reg_r_9[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_8 = result_reg_r_9[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_9 = result_reg_r_9[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_10 = result_reg_r_9[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_11 = result_reg_r_9[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_12 = result_reg_r_9[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_13 = result_reg_r_9[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_14 = result_reg_r_9[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_15 = result_reg_r_9[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_16 = result_reg_r_9[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_17 = result_reg_r_9[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_18 = result_reg_r_9[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_19 = result_reg_r_9[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_20 = result_reg_r_9[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_21 = result_reg_r_9[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_22 = result_reg_r_9[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_23 = result_reg_r_9[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_24 = result_reg_r_9[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_25 = result_reg_r_9[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_26 = result_reg_r_9[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_27 = result_reg_r_9[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_28 = result_reg_r_9[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_29 = result_reg_r_9[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_30 = result_reg_r_9[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_31 = result_reg_r_9[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_32 = result_reg_r_9[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_33 = result_reg_r_9[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_34 = result_reg_r_9[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_35 = result_reg_r_9[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_36 = result_reg_r_9[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_37 = result_reg_r_9[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_38 = result_reg_r_9[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_39 = result_reg_r_9[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_40 = result_reg_r_9[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_41 = result_reg_r_9[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_42 = result_reg_r_9[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_43 = result_reg_r_9[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_44 = result_reg_r_9[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_45 = result_reg_r_9[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_46 = result_reg_r_9[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_47 = result_reg_r_9[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_48 = result_reg_r_9[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_49 = result_reg_r_9[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_50 = result_reg_r_9[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_51 = result_reg_r_9[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_52 = result_reg_r_9[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_53 = result_reg_r_9[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_54 = result_reg_r_9[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_55 = result_reg_r_9[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_56 = result_reg_r_9[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_57 = result_reg_r_9[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_58 = result_reg_r_9[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_59 = result_reg_r_9[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_60 = result_reg_r_9[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_61 = result_reg_r_9[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_62 = result_reg_r_9[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_63 = result_reg_r_9[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_64 = result_reg_r_9[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_65 = result_reg_r_9[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_66 = result_reg_r_9[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_67 = result_reg_r_9[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_68 = result_reg_r_9[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_69 = result_reg_r_9[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_70 = result_reg_r_9[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_71 = result_reg_r_9[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_72 = result_reg_r_9[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_73 = result_reg_r_9[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_74 = result_reg_r_9[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_75 = result_reg_r_9[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_76 = result_reg_r_9[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_77 = result_reg_r_9[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_78 = result_reg_r_9[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_79 = result_reg_r_9[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_80 = result_reg_r_9[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_81 = result_reg_r_9[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_82 = result_reg_r_9[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_83 = result_reg_r_9[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_84 = result_reg_r_9[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_86 = result_reg_r_9[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_87 = result_reg_r_9[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_88 = result_reg_r_9[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_89 = result_reg_r_9[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_90 = result_reg_r_9[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_91 = result_reg_r_9[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_92 = result_reg_r_9[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_93 = result_reg_r_9[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_94 = result_reg_r_9[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_95 = result_reg_r_9[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_96 = result_reg_r_9[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_97 = result_reg_r_9[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_98 = result_reg_r_9[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_99 = result_reg_r_9[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_100 = result_reg_r_9[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_101 = result_reg_r_9[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_102 = result_reg_r_9[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_103 = result_reg_r_9[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_104 = result_reg_r_9[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_19_105 = result_reg_r_9[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_10_hi_hi_hi_lo = {wire_res_19_98,wire_res_19_97,wire_res_19_96,wire_res_19_95,wire_res_19_94,
    wire_res_19_93,wire_res_19_92}; // @[BinaryDesigns2.scala 231:46]
  wire [190:0] _T_11276 = {b_aux_reg_r_9, 85'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [190:0] _GEN_1281 = {{85'd0}, a_aux_reg_r_9}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_19_85 = _GEN_1281 >= _T_11276; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_10_hi_hi_lo_lo = {wire_res_19_84,wire_res_19_83,wire_res_19_82,wire_res_19_81,wire_res_19_80,
    wire_res_19_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_10_hi_hi_lo = {wire_res_19_91,wire_res_19_90,wire_res_19_89,wire_res_19_88,wire_res_19_87,
    wire_res_19_86,wire_res_19_85,result_reg_w_10_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_10_hi_lo_hi_lo = {wire_res_19_71,wire_res_19_70,wire_res_19_69,wire_res_19_68,wire_res_19_67,
    wire_res_19_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_10_hi_lo_lo_lo = {wire_res_19_58,wire_res_19_57,wire_res_19_56,wire_res_19_55,wire_res_19_54,
    wire_res_19_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_10_hi_lo_lo = {wire_res_19_65,wire_res_19_64,wire_res_19_63,wire_res_19_62,wire_res_19_61,
    wire_res_19_60,wire_res_19_59,result_reg_w_10_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_10_hi_lo = {wire_res_19_78,wire_res_19_77,wire_res_19_76,wire_res_19_75,wire_res_19_74,
    wire_res_19_73,wire_res_19_72,result_reg_w_10_hi_lo_hi_lo,result_reg_w_10_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_10_hi = {wire_res_19_105,wire_res_19_104,wire_res_19_103,wire_res_19_102,wire_res_19_101,
    wire_res_19_100,wire_res_19_99,result_reg_w_10_hi_hi_hi_lo,result_reg_w_10_hi_hi_lo,result_reg_w_10_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_10_lo_hi_hi_lo = {wire_res_19_45,wire_res_19_44,wire_res_19_43,wire_res_19_42,wire_res_19_41,
    wire_res_19_40,wire_res_19_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_10_lo_hi_lo_lo = {wire_res_19_31,wire_res_19_30,wire_res_19_29,wire_res_19_28,wire_res_19_27,
    wire_res_19_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_10_lo_hi_lo = {wire_res_19_38,wire_res_19_37,wire_res_19_36,wire_res_19_35,wire_res_19_34,
    wire_res_19_33,wire_res_19_32,result_reg_w_10_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_10_lo_lo_hi_lo = {wire_res_19_18,wire_res_19_17,wire_res_19_16,wire_res_19_15,wire_res_19_14,
    wire_res_19_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_10_lo_lo_lo_lo = {wire_res_19_5,wire_res_19_4,wire_res_19_3,wire_res_19_2,wire_res_19_1,
    wire_res_19_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_10_lo_lo_lo = {wire_res_19_12,wire_res_19_11,wire_res_19_10,wire_res_19_9,wire_res_19_8,
    wire_res_19_7,wire_res_19_6,result_reg_w_10_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_10_lo_lo = {wire_res_19_25,wire_res_19_24,wire_res_19_23,wire_res_19_22,wire_res_19_21,
    wire_res_19_20,wire_res_19_19,result_reg_w_10_lo_lo_hi_lo,result_reg_w_10_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_10_lo = {wire_res_19_52,wire_res_19_51,wire_res_19_50,wire_res_19_49,wire_res_19_48,
    wire_res_19_47,wire_res_19_46,result_reg_w_10_lo_hi_hi_lo,result_reg_w_10_lo_hi_lo,result_reg_w_10_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_10 = {result_reg_w_10_hi,result_reg_w_10_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_20_0 = result_reg_w_10[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_1 = result_reg_w_10[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_2 = result_reg_w_10[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_3 = result_reg_w_10[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_4 = result_reg_w_10[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_5 = result_reg_w_10[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_6 = result_reg_w_10[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_7 = result_reg_w_10[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_8 = result_reg_w_10[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_9 = result_reg_w_10[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_10 = result_reg_w_10[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_11 = result_reg_w_10[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_12 = result_reg_w_10[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_13 = result_reg_w_10[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_14 = result_reg_w_10[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_15 = result_reg_w_10[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_16 = result_reg_w_10[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_17 = result_reg_w_10[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_18 = result_reg_w_10[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_19 = result_reg_w_10[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_20 = result_reg_w_10[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_21 = result_reg_w_10[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_22 = result_reg_w_10[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_23 = result_reg_w_10[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_24 = result_reg_w_10[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_25 = result_reg_w_10[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_26 = result_reg_w_10[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_27 = result_reg_w_10[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_28 = result_reg_w_10[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_29 = result_reg_w_10[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_30 = result_reg_w_10[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_31 = result_reg_w_10[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_32 = result_reg_w_10[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_33 = result_reg_w_10[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_34 = result_reg_w_10[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_35 = result_reg_w_10[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_36 = result_reg_w_10[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_37 = result_reg_w_10[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_38 = result_reg_w_10[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_39 = result_reg_w_10[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_40 = result_reg_w_10[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_41 = result_reg_w_10[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_42 = result_reg_w_10[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_43 = result_reg_w_10[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_44 = result_reg_w_10[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_45 = result_reg_w_10[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_46 = result_reg_w_10[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_47 = result_reg_w_10[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_48 = result_reg_w_10[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_49 = result_reg_w_10[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_50 = result_reg_w_10[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_51 = result_reg_w_10[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_52 = result_reg_w_10[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_53 = result_reg_w_10[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_54 = result_reg_w_10[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_55 = result_reg_w_10[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_56 = result_reg_w_10[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_57 = result_reg_w_10[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_58 = result_reg_w_10[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_59 = result_reg_w_10[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_60 = result_reg_w_10[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_61 = result_reg_w_10[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_62 = result_reg_w_10[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_63 = result_reg_w_10[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_64 = result_reg_w_10[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_65 = result_reg_w_10[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_66 = result_reg_w_10[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_67 = result_reg_w_10[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_68 = result_reg_w_10[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_69 = result_reg_w_10[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_70 = result_reg_w_10[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_71 = result_reg_w_10[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_72 = result_reg_w_10[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_73 = result_reg_w_10[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_74 = result_reg_w_10[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_75 = result_reg_w_10[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_76 = result_reg_w_10[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_77 = result_reg_w_10[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_78 = result_reg_w_10[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_79 = result_reg_w_10[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_80 = result_reg_w_10[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_81 = result_reg_w_10[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_82 = result_reg_w_10[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_83 = result_reg_w_10[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_85 = result_reg_w_10[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_86 = result_reg_w_10[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_87 = result_reg_w_10[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_88 = result_reg_w_10[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_89 = result_reg_w_10[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_90 = result_reg_w_10[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_91 = result_reg_w_10[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_92 = result_reg_w_10[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_93 = result_reg_w_10[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_94 = result_reg_w_10[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_95 = result_reg_w_10[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_96 = result_reg_w_10[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_97 = result_reg_w_10[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_98 = result_reg_w_10[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_99 = result_reg_w_10[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_100 = result_reg_w_10[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_101 = result_reg_w_10[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_102 = result_reg_w_10[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_103 = result_reg_w_10[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_104 = result_reg_w_10[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_20_105 = result_reg_w_10[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_0 = result_reg_r_10[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_1 = result_reg_r_10[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_2 = result_reg_r_10[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_3 = result_reg_r_10[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_4 = result_reg_r_10[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_5 = result_reg_r_10[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_6 = result_reg_r_10[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_7 = result_reg_r_10[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_8 = result_reg_r_10[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_9 = result_reg_r_10[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_10 = result_reg_r_10[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_11 = result_reg_r_10[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_12 = result_reg_r_10[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_13 = result_reg_r_10[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_14 = result_reg_r_10[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_15 = result_reg_r_10[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_16 = result_reg_r_10[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_17 = result_reg_r_10[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_18 = result_reg_r_10[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_19 = result_reg_r_10[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_20 = result_reg_r_10[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_21 = result_reg_r_10[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_22 = result_reg_r_10[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_23 = result_reg_r_10[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_24 = result_reg_r_10[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_25 = result_reg_r_10[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_26 = result_reg_r_10[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_27 = result_reg_r_10[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_28 = result_reg_r_10[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_29 = result_reg_r_10[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_30 = result_reg_r_10[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_31 = result_reg_r_10[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_32 = result_reg_r_10[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_33 = result_reg_r_10[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_34 = result_reg_r_10[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_35 = result_reg_r_10[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_36 = result_reg_r_10[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_37 = result_reg_r_10[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_38 = result_reg_r_10[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_39 = result_reg_r_10[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_40 = result_reg_r_10[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_41 = result_reg_r_10[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_42 = result_reg_r_10[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_43 = result_reg_r_10[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_44 = result_reg_r_10[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_45 = result_reg_r_10[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_46 = result_reg_r_10[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_47 = result_reg_r_10[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_48 = result_reg_r_10[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_49 = result_reg_r_10[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_50 = result_reg_r_10[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_51 = result_reg_r_10[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_52 = result_reg_r_10[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_53 = result_reg_r_10[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_54 = result_reg_r_10[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_55 = result_reg_r_10[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_56 = result_reg_r_10[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_57 = result_reg_r_10[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_58 = result_reg_r_10[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_59 = result_reg_r_10[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_60 = result_reg_r_10[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_61 = result_reg_r_10[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_62 = result_reg_r_10[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_63 = result_reg_r_10[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_64 = result_reg_r_10[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_65 = result_reg_r_10[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_66 = result_reg_r_10[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_67 = result_reg_r_10[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_68 = result_reg_r_10[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_69 = result_reg_r_10[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_70 = result_reg_r_10[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_71 = result_reg_r_10[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_72 = result_reg_r_10[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_73 = result_reg_r_10[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_74 = result_reg_r_10[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_75 = result_reg_r_10[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_76 = result_reg_r_10[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_77 = result_reg_r_10[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_78 = result_reg_r_10[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_79 = result_reg_r_10[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_80 = result_reg_r_10[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_81 = result_reg_r_10[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_82 = result_reg_r_10[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_84 = result_reg_r_10[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_85 = result_reg_r_10[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_86 = result_reg_r_10[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_87 = result_reg_r_10[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_88 = result_reg_r_10[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_89 = result_reg_r_10[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_90 = result_reg_r_10[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_91 = result_reg_r_10[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_92 = result_reg_r_10[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_93 = result_reg_r_10[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_94 = result_reg_r_10[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_95 = result_reg_r_10[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_96 = result_reg_r_10[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_97 = result_reg_r_10[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_98 = result_reg_r_10[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_99 = result_reg_r_10[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_100 = result_reg_r_10[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_101 = result_reg_r_10[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_102 = result_reg_r_10[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_103 = result_reg_r_10[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_104 = result_reg_r_10[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_21_105 = result_reg_r_10[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_11_hi_hi_hi_lo = {wire_res_21_98,wire_res_21_97,wire_res_21_96,wire_res_21_95,wire_res_21_94,
    wire_res_21_93,wire_res_21_92}; // @[BinaryDesigns2.scala 231:46]
  wire [188:0] _T_11280 = {b_aux_reg_r_10, 83'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [188:0] _GEN_1282 = {{83'd0}, a_aux_reg_r_10}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_21_83 = _GEN_1282 >= _T_11280; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_11_hi_hi_lo_lo = {wire_res_21_84,wire_res_21_83,wire_res_21_82,wire_res_21_81,wire_res_21_80,
    wire_res_21_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_11_hi_hi_lo = {wire_res_21_91,wire_res_21_90,wire_res_21_89,wire_res_21_88,wire_res_21_87,
    wire_res_21_86,wire_res_21_85,result_reg_w_11_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_11_hi_lo_hi_lo = {wire_res_21_71,wire_res_21_70,wire_res_21_69,wire_res_21_68,wire_res_21_67,
    wire_res_21_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_11_hi_lo_lo_lo = {wire_res_21_58,wire_res_21_57,wire_res_21_56,wire_res_21_55,wire_res_21_54,
    wire_res_21_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_11_hi_lo_lo = {wire_res_21_65,wire_res_21_64,wire_res_21_63,wire_res_21_62,wire_res_21_61,
    wire_res_21_60,wire_res_21_59,result_reg_w_11_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_11_hi_lo = {wire_res_21_78,wire_res_21_77,wire_res_21_76,wire_res_21_75,wire_res_21_74,
    wire_res_21_73,wire_res_21_72,result_reg_w_11_hi_lo_hi_lo,result_reg_w_11_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_11_hi = {wire_res_21_105,wire_res_21_104,wire_res_21_103,wire_res_21_102,wire_res_21_101,
    wire_res_21_100,wire_res_21_99,result_reg_w_11_hi_hi_hi_lo,result_reg_w_11_hi_hi_lo,result_reg_w_11_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_11_lo_hi_hi_lo = {wire_res_21_45,wire_res_21_44,wire_res_21_43,wire_res_21_42,wire_res_21_41,
    wire_res_21_40,wire_res_21_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_11_lo_hi_lo_lo = {wire_res_21_31,wire_res_21_30,wire_res_21_29,wire_res_21_28,wire_res_21_27,
    wire_res_21_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_11_lo_hi_lo = {wire_res_21_38,wire_res_21_37,wire_res_21_36,wire_res_21_35,wire_res_21_34,
    wire_res_21_33,wire_res_21_32,result_reg_w_11_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_11_lo_lo_hi_lo = {wire_res_21_18,wire_res_21_17,wire_res_21_16,wire_res_21_15,wire_res_21_14,
    wire_res_21_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_11_lo_lo_lo_lo = {wire_res_21_5,wire_res_21_4,wire_res_21_3,wire_res_21_2,wire_res_21_1,
    wire_res_21_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_11_lo_lo_lo = {wire_res_21_12,wire_res_21_11,wire_res_21_10,wire_res_21_9,wire_res_21_8,
    wire_res_21_7,wire_res_21_6,result_reg_w_11_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_11_lo_lo = {wire_res_21_25,wire_res_21_24,wire_res_21_23,wire_res_21_22,wire_res_21_21,
    wire_res_21_20,wire_res_21_19,result_reg_w_11_lo_lo_hi_lo,result_reg_w_11_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_11_lo = {wire_res_21_52,wire_res_21_51,wire_res_21_50,wire_res_21_49,wire_res_21_48,
    wire_res_21_47,wire_res_21_46,result_reg_w_11_lo_hi_hi_lo,result_reg_w_11_lo_hi_lo,result_reg_w_11_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_11 = {result_reg_w_11_hi,result_reg_w_11_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_22_0 = result_reg_w_11[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_1 = result_reg_w_11[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_2 = result_reg_w_11[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_3 = result_reg_w_11[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_4 = result_reg_w_11[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_5 = result_reg_w_11[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_6 = result_reg_w_11[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_7 = result_reg_w_11[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_8 = result_reg_w_11[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_9 = result_reg_w_11[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_10 = result_reg_w_11[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_11 = result_reg_w_11[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_12 = result_reg_w_11[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_13 = result_reg_w_11[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_14 = result_reg_w_11[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_15 = result_reg_w_11[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_16 = result_reg_w_11[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_17 = result_reg_w_11[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_18 = result_reg_w_11[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_19 = result_reg_w_11[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_20 = result_reg_w_11[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_21 = result_reg_w_11[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_22 = result_reg_w_11[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_23 = result_reg_w_11[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_24 = result_reg_w_11[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_25 = result_reg_w_11[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_26 = result_reg_w_11[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_27 = result_reg_w_11[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_28 = result_reg_w_11[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_29 = result_reg_w_11[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_30 = result_reg_w_11[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_31 = result_reg_w_11[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_32 = result_reg_w_11[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_33 = result_reg_w_11[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_34 = result_reg_w_11[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_35 = result_reg_w_11[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_36 = result_reg_w_11[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_37 = result_reg_w_11[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_38 = result_reg_w_11[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_39 = result_reg_w_11[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_40 = result_reg_w_11[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_41 = result_reg_w_11[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_42 = result_reg_w_11[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_43 = result_reg_w_11[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_44 = result_reg_w_11[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_45 = result_reg_w_11[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_46 = result_reg_w_11[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_47 = result_reg_w_11[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_48 = result_reg_w_11[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_49 = result_reg_w_11[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_50 = result_reg_w_11[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_51 = result_reg_w_11[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_52 = result_reg_w_11[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_53 = result_reg_w_11[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_54 = result_reg_w_11[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_55 = result_reg_w_11[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_56 = result_reg_w_11[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_57 = result_reg_w_11[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_58 = result_reg_w_11[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_59 = result_reg_w_11[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_60 = result_reg_w_11[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_61 = result_reg_w_11[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_62 = result_reg_w_11[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_63 = result_reg_w_11[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_64 = result_reg_w_11[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_65 = result_reg_w_11[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_66 = result_reg_w_11[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_67 = result_reg_w_11[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_68 = result_reg_w_11[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_69 = result_reg_w_11[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_70 = result_reg_w_11[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_71 = result_reg_w_11[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_72 = result_reg_w_11[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_73 = result_reg_w_11[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_74 = result_reg_w_11[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_75 = result_reg_w_11[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_76 = result_reg_w_11[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_77 = result_reg_w_11[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_78 = result_reg_w_11[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_79 = result_reg_w_11[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_80 = result_reg_w_11[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_81 = result_reg_w_11[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_83 = result_reg_w_11[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_84 = result_reg_w_11[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_85 = result_reg_w_11[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_86 = result_reg_w_11[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_87 = result_reg_w_11[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_88 = result_reg_w_11[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_89 = result_reg_w_11[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_90 = result_reg_w_11[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_91 = result_reg_w_11[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_92 = result_reg_w_11[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_93 = result_reg_w_11[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_94 = result_reg_w_11[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_95 = result_reg_w_11[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_96 = result_reg_w_11[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_97 = result_reg_w_11[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_98 = result_reg_w_11[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_99 = result_reg_w_11[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_100 = result_reg_w_11[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_101 = result_reg_w_11[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_102 = result_reg_w_11[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_103 = result_reg_w_11[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_104 = result_reg_w_11[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_22_105 = result_reg_w_11[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_0 = result_reg_r_11[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_1 = result_reg_r_11[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_2 = result_reg_r_11[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_3 = result_reg_r_11[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_4 = result_reg_r_11[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_5 = result_reg_r_11[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_6 = result_reg_r_11[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_7 = result_reg_r_11[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_8 = result_reg_r_11[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_9 = result_reg_r_11[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_10 = result_reg_r_11[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_11 = result_reg_r_11[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_12 = result_reg_r_11[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_13 = result_reg_r_11[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_14 = result_reg_r_11[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_15 = result_reg_r_11[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_16 = result_reg_r_11[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_17 = result_reg_r_11[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_18 = result_reg_r_11[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_19 = result_reg_r_11[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_20 = result_reg_r_11[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_21 = result_reg_r_11[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_22 = result_reg_r_11[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_23 = result_reg_r_11[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_24 = result_reg_r_11[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_25 = result_reg_r_11[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_26 = result_reg_r_11[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_27 = result_reg_r_11[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_28 = result_reg_r_11[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_29 = result_reg_r_11[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_30 = result_reg_r_11[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_31 = result_reg_r_11[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_32 = result_reg_r_11[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_33 = result_reg_r_11[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_34 = result_reg_r_11[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_35 = result_reg_r_11[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_36 = result_reg_r_11[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_37 = result_reg_r_11[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_38 = result_reg_r_11[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_39 = result_reg_r_11[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_40 = result_reg_r_11[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_41 = result_reg_r_11[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_42 = result_reg_r_11[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_43 = result_reg_r_11[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_44 = result_reg_r_11[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_45 = result_reg_r_11[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_46 = result_reg_r_11[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_47 = result_reg_r_11[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_48 = result_reg_r_11[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_49 = result_reg_r_11[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_50 = result_reg_r_11[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_51 = result_reg_r_11[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_52 = result_reg_r_11[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_53 = result_reg_r_11[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_54 = result_reg_r_11[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_55 = result_reg_r_11[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_56 = result_reg_r_11[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_57 = result_reg_r_11[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_58 = result_reg_r_11[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_59 = result_reg_r_11[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_60 = result_reg_r_11[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_61 = result_reg_r_11[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_62 = result_reg_r_11[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_63 = result_reg_r_11[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_64 = result_reg_r_11[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_65 = result_reg_r_11[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_66 = result_reg_r_11[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_67 = result_reg_r_11[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_68 = result_reg_r_11[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_69 = result_reg_r_11[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_70 = result_reg_r_11[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_71 = result_reg_r_11[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_72 = result_reg_r_11[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_73 = result_reg_r_11[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_74 = result_reg_r_11[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_75 = result_reg_r_11[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_76 = result_reg_r_11[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_77 = result_reg_r_11[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_78 = result_reg_r_11[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_79 = result_reg_r_11[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_80 = result_reg_r_11[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_82 = result_reg_r_11[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_83 = result_reg_r_11[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_84 = result_reg_r_11[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_85 = result_reg_r_11[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_86 = result_reg_r_11[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_87 = result_reg_r_11[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_88 = result_reg_r_11[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_89 = result_reg_r_11[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_90 = result_reg_r_11[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_91 = result_reg_r_11[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_92 = result_reg_r_11[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_93 = result_reg_r_11[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_94 = result_reg_r_11[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_95 = result_reg_r_11[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_96 = result_reg_r_11[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_97 = result_reg_r_11[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_98 = result_reg_r_11[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_99 = result_reg_r_11[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_100 = result_reg_r_11[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_101 = result_reg_r_11[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_102 = result_reg_r_11[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_103 = result_reg_r_11[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_104 = result_reg_r_11[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_23_105 = result_reg_r_11[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_12_hi_hi_hi_lo = {wire_res_23_98,wire_res_23_97,wire_res_23_96,wire_res_23_95,wire_res_23_94,
    wire_res_23_93,wire_res_23_92}; // @[BinaryDesigns2.scala 231:46]
  wire [186:0] _T_11284 = {b_aux_reg_r_11, 81'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [186:0] _GEN_1283 = {{81'd0}, a_aux_reg_r_11}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_23_81 = _GEN_1283 >= _T_11284; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_12_hi_hi_lo_lo = {wire_res_23_84,wire_res_23_83,wire_res_23_82,wire_res_23_81,wire_res_23_80,
    wire_res_23_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_12_hi_hi_lo = {wire_res_23_91,wire_res_23_90,wire_res_23_89,wire_res_23_88,wire_res_23_87,
    wire_res_23_86,wire_res_23_85,result_reg_w_12_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_12_hi_lo_hi_lo = {wire_res_23_71,wire_res_23_70,wire_res_23_69,wire_res_23_68,wire_res_23_67,
    wire_res_23_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_12_hi_lo_lo_lo = {wire_res_23_58,wire_res_23_57,wire_res_23_56,wire_res_23_55,wire_res_23_54,
    wire_res_23_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_12_hi_lo_lo = {wire_res_23_65,wire_res_23_64,wire_res_23_63,wire_res_23_62,wire_res_23_61,
    wire_res_23_60,wire_res_23_59,result_reg_w_12_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_12_hi_lo = {wire_res_23_78,wire_res_23_77,wire_res_23_76,wire_res_23_75,wire_res_23_74,
    wire_res_23_73,wire_res_23_72,result_reg_w_12_hi_lo_hi_lo,result_reg_w_12_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_12_hi = {wire_res_23_105,wire_res_23_104,wire_res_23_103,wire_res_23_102,wire_res_23_101,
    wire_res_23_100,wire_res_23_99,result_reg_w_12_hi_hi_hi_lo,result_reg_w_12_hi_hi_lo,result_reg_w_12_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_12_lo_hi_hi_lo = {wire_res_23_45,wire_res_23_44,wire_res_23_43,wire_res_23_42,wire_res_23_41,
    wire_res_23_40,wire_res_23_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_12_lo_hi_lo_lo = {wire_res_23_31,wire_res_23_30,wire_res_23_29,wire_res_23_28,wire_res_23_27,
    wire_res_23_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_12_lo_hi_lo = {wire_res_23_38,wire_res_23_37,wire_res_23_36,wire_res_23_35,wire_res_23_34,
    wire_res_23_33,wire_res_23_32,result_reg_w_12_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_12_lo_lo_hi_lo = {wire_res_23_18,wire_res_23_17,wire_res_23_16,wire_res_23_15,wire_res_23_14,
    wire_res_23_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_12_lo_lo_lo_lo = {wire_res_23_5,wire_res_23_4,wire_res_23_3,wire_res_23_2,wire_res_23_1,
    wire_res_23_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_12_lo_lo_lo = {wire_res_23_12,wire_res_23_11,wire_res_23_10,wire_res_23_9,wire_res_23_8,
    wire_res_23_7,wire_res_23_6,result_reg_w_12_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_12_lo_lo = {wire_res_23_25,wire_res_23_24,wire_res_23_23,wire_res_23_22,wire_res_23_21,
    wire_res_23_20,wire_res_23_19,result_reg_w_12_lo_lo_hi_lo,result_reg_w_12_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_12_lo = {wire_res_23_52,wire_res_23_51,wire_res_23_50,wire_res_23_49,wire_res_23_48,
    wire_res_23_47,wire_res_23_46,result_reg_w_12_lo_hi_hi_lo,result_reg_w_12_lo_hi_lo,result_reg_w_12_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_12 = {result_reg_w_12_hi,result_reg_w_12_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_24_0 = result_reg_w_12[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_1 = result_reg_w_12[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_2 = result_reg_w_12[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_3 = result_reg_w_12[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_4 = result_reg_w_12[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_5 = result_reg_w_12[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_6 = result_reg_w_12[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_7 = result_reg_w_12[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_8 = result_reg_w_12[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_9 = result_reg_w_12[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_10 = result_reg_w_12[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_11 = result_reg_w_12[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_12 = result_reg_w_12[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_13 = result_reg_w_12[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_14 = result_reg_w_12[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_15 = result_reg_w_12[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_16 = result_reg_w_12[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_17 = result_reg_w_12[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_18 = result_reg_w_12[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_19 = result_reg_w_12[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_20 = result_reg_w_12[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_21 = result_reg_w_12[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_22 = result_reg_w_12[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_23 = result_reg_w_12[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_24 = result_reg_w_12[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_25 = result_reg_w_12[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_26 = result_reg_w_12[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_27 = result_reg_w_12[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_28 = result_reg_w_12[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_29 = result_reg_w_12[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_30 = result_reg_w_12[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_31 = result_reg_w_12[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_32 = result_reg_w_12[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_33 = result_reg_w_12[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_34 = result_reg_w_12[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_35 = result_reg_w_12[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_36 = result_reg_w_12[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_37 = result_reg_w_12[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_38 = result_reg_w_12[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_39 = result_reg_w_12[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_40 = result_reg_w_12[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_41 = result_reg_w_12[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_42 = result_reg_w_12[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_43 = result_reg_w_12[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_44 = result_reg_w_12[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_45 = result_reg_w_12[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_46 = result_reg_w_12[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_47 = result_reg_w_12[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_48 = result_reg_w_12[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_49 = result_reg_w_12[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_50 = result_reg_w_12[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_51 = result_reg_w_12[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_52 = result_reg_w_12[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_53 = result_reg_w_12[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_54 = result_reg_w_12[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_55 = result_reg_w_12[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_56 = result_reg_w_12[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_57 = result_reg_w_12[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_58 = result_reg_w_12[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_59 = result_reg_w_12[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_60 = result_reg_w_12[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_61 = result_reg_w_12[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_62 = result_reg_w_12[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_63 = result_reg_w_12[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_64 = result_reg_w_12[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_65 = result_reg_w_12[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_66 = result_reg_w_12[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_67 = result_reg_w_12[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_68 = result_reg_w_12[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_69 = result_reg_w_12[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_70 = result_reg_w_12[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_71 = result_reg_w_12[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_72 = result_reg_w_12[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_73 = result_reg_w_12[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_74 = result_reg_w_12[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_75 = result_reg_w_12[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_76 = result_reg_w_12[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_77 = result_reg_w_12[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_78 = result_reg_w_12[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_79 = result_reg_w_12[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_81 = result_reg_w_12[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_82 = result_reg_w_12[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_83 = result_reg_w_12[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_84 = result_reg_w_12[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_85 = result_reg_w_12[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_86 = result_reg_w_12[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_87 = result_reg_w_12[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_88 = result_reg_w_12[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_89 = result_reg_w_12[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_90 = result_reg_w_12[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_91 = result_reg_w_12[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_92 = result_reg_w_12[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_93 = result_reg_w_12[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_94 = result_reg_w_12[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_95 = result_reg_w_12[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_96 = result_reg_w_12[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_97 = result_reg_w_12[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_98 = result_reg_w_12[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_99 = result_reg_w_12[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_100 = result_reg_w_12[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_101 = result_reg_w_12[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_102 = result_reg_w_12[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_103 = result_reg_w_12[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_104 = result_reg_w_12[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_24_105 = result_reg_w_12[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_0 = result_reg_r_12[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_1 = result_reg_r_12[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_2 = result_reg_r_12[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_3 = result_reg_r_12[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_4 = result_reg_r_12[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_5 = result_reg_r_12[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_6 = result_reg_r_12[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_7 = result_reg_r_12[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_8 = result_reg_r_12[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_9 = result_reg_r_12[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_10 = result_reg_r_12[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_11 = result_reg_r_12[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_12 = result_reg_r_12[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_13 = result_reg_r_12[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_14 = result_reg_r_12[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_15 = result_reg_r_12[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_16 = result_reg_r_12[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_17 = result_reg_r_12[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_18 = result_reg_r_12[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_19 = result_reg_r_12[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_20 = result_reg_r_12[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_21 = result_reg_r_12[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_22 = result_reg_r_12[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_23 = result_reg_r_12[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_24 = result_reg_r_12[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_25 = result_reg_r_12[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_26 = result_reg_r_12[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_27 = result_reg_r_12[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_28 = result_reg_r_12[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_29 = result_reg_r_12[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_30 = result_reg_r_12[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_31 = result_reg_r_12[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_32 = result_reg_r_12[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_33 = result_reg_r_12[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_34 = result_reg_r_12[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_35 = result_reg_r_12[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_36 = result_reg_r_12[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_37 = result_reg_r_12[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_38 = result_reg_r_12[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_39 = result_reg_r_12[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_40 = result_reg_r_12[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_41 = result_reg_r_12[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_42 = result_reg_r_12[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_43 = result_reg_r_12[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_44 = result_reg_r_12[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_45 = result_reg_r_12[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_46 = result_reg_r_12[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_47 = result_reg_r_12[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_48 = result_reg_r_12[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_49 = result_reg_r_12[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_50 = result_reg_r_12[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_51 = result_reg_r_12[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_52 = result_reg_r_12[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_53 = result_reg_r_12[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_54 = result_reg_r_12[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_55 = result_reg_r_12[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_56 = result_reg_r_12[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_57 = result_reg_r_12[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_58 = result_reg_r_12[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_59 = result_reg_r_12[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_60 = result_reg_r_12[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_61 = result_reg_r_12[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_62 = result_reg_r_12[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_63 = result_reg_r_12[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_64 = result_reg_r_12[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_65 = result_reg_r_12[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_66 = result_reg_r_12[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_67 = result_reg_r_12[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_68 = result_reg_r_12[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_69 = result_reg_r_12[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_70 = result_reg_r_12[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_71 = result_reg_r_12[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_72 = result_reg_r_12[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_73 = result_reg_r_12[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_74 = result_reg_r_12[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_75 = result_reg_r_12[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_76 = result_reg_r_12[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_77 = result_reg_r_12[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_78 = result_reg_r_12[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_80 = result_reg_r_12[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_81 = result_reg_r_12[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_82 = result_reg_r_12[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_83 = result_reg_r_12[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_84 = result_reg_r_12[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_85 = result_reg_r_12[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_86 = result_reg_r_12[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_87 = result_reg_r_12[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_88 = result_reg_r_12[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_89 = result_reg_r_12[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_90 = result_reg_r_12[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_91 = result_reg_r_12[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_92 = result_reg_r_12[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_93 = result_reg_r_12[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_94 = result_reg_r_12[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_95 = result_reg_r_12[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_96 = result_reg_r_12[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_97 = result_reg_r_12[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_98 = result_reg_r_12[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_99 = result_reg_r_12[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_100 = result_reg_r_12[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_101 = result_reg_r_12[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_102 = result_reg_r_12[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_103 = result_reg_r_12[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_104 = result_reg_r_12[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_25_105 = result_reg_r_12[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_13_hi_hi_hi_lo = {wire_res_25_98,wire_res_25_97,wire_res_25_96,wire_res_25_95,wire_res_25_94,
    wire_res_25_93,wire_res_25_92}; // @[BinaryDesigns2.scala 231:46]
  wire [184:0] _T_11288 = {b_aux_reg_r_12, 79'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [184:0] _GEN_1284 = {{79'd0}, a_aux_reg_r_12}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_25_79 = _GEN_1284 >= _T_11288; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_13_hi_hi_lo_lo = {wire_res_25_84,wire_res_25_83,wire_res_25_82,wire_res_25_81,wire_res_25_80,
    wire_res_25_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_13_hi_hi_lo = {wire_res_25_91,wire_res_25_90,wire_res_25_89,wire_res_25_88,wire_res_25_87,
    wire_res_25_86,wire_res_25_85,result_reg_w_13_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_13_hi_lo_hi_lo = {wire_res_25_71,wire_res_25_70,wire_res_25_69,wire_res_25_68,wire_res_25_67,
    wire_res_25_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_13_hi_lo_lo_lo = {wire_res_25_58,wire_res_25_57,wire_res_25_56,wire_res_25_55,wire_res_25_54,
    wire_res_25_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_13_hi_lo_lo = {wire_res_25_65,wire_res_25_64,wire_res_25_63,wire_res_25_62,wire_res_25_61,
    wire_res_25_60,wire_res_25_59,result_reg_w_13_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_13_hi_lo = {wire_res_25_78,wire_res_25_77,wire_res_25_76,wire_res_25_75,wire_res_25_74,
    wire_res_25_73,wire_res_25_72,result_reg_w_13_hi_lo_hi_lo,result_reg_w_13_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_13_hi = {wire_res_25_105,wire_res_25_104,wire_res_25_103,wire_res_25_102,wire_res_25_101,
    wire_res_25_100,wire_res_25_99,result_reg_w_13_hi_hi_hi_lo,result_reg_w_13_hi_hi_lo,result_reg_w_13_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_13_lo_hi_hi_lo = {wire_res_25_45,wire_res_25_44,wire_res_25_43,wire_res_25_42,wire_res_25_41,
    wire_res_25_40,wire_res_25_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_13_lo_hi_lo_lo = {wire_res_25_31,wire_res_25_30,wire_res_25_29,wire_res_25_28,wire_res_25_27,
    wire_res_25_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_13_lo_hi_lo = {wire_res_25_38,wire_res_25_37,wire_res_25_36,wire_res_25_35,wire_res_25_34,
    wire_res_25_33,wire_res_25_32,result_reg_w_13_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_13_lo_lo_hi_lo = {wire_res_25_18,wire_res_25_17,wire_res_25_16,wire_res_25_15,wire_res_25_14,
    wire_res_25_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_13_lo_lo_lo_lo = {wire_res_25_5,wire_res_25_4,wire_res_25_3,wire_res_25_2,wire_res_25_1,
    wire_res_25_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_13_lo_lo_lo = {wire_res_25_12,wire_res_25_11,wire_res_25_10,wire_res_25_9,wire_res_25_8,
    wire_res_25_7,wire_res_25_6,result_reg_w_13_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_13_lo_lo = {wire_res_25_25,wire_res_25_24,wire_res_25_23,wire_res_25_22,wire_res_25_21,
    wire_res_25_20,wire_res_25_19,result_reg_w_13_lo_lo_hi_lo,result_reg_w_13_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_13_lo = {wire_res_25_52,wire_res_25_51,wire_res_25_50,wire_res_25_49,wire_res_25_48,
    wire_res_25_47,wire_res_25_46,result_reg_w_13_lo_hi_hi_lo,result_reg_w_13_lo_hi_lo,result_reg_w_13_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_13 = {result_reg_w_13_hi,result_reg_w_13_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_26_0 = result_reg_w_13[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_1 = result_reg_w_13[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_2 = result_reg_w_13[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_3 = result_reg_w_13[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_4 = result_reg_w_13[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_5 = result_reg_w_13[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_6 = result_reg_w_13[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_7 = result_reg_w_13[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_8 = result_reg_w_13[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_9 = result_reg_w_13[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_10 = result_reg_w_13[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_11 = result_reg_w_13[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_12 = result_reg_w_13[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_13 = result_reg_w_13[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_14 = result_reg_w_13[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_15 = result_reg_w_13[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_16 = result_reg_w_13[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_17 = result_reg_w_13[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_18 = result_reg_w_13[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_19 = result_reg_w_13[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_20 = result_reg_w_13[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_21 = result_reg_w_13[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_22 = result_reg_w_13[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_23 = result_reg_w_13[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_24 = result_reg_w_13[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_25 = result_reg_w_13[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_26 = result_reg_w_13[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_27 = result_reg_w_13[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_28 = result_reg_w_13[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_29 = result_reg_w_13[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_30 = result_reg_w_13[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_31 = result_reg_w_13[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_32 = result_reg_w_13[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_33 = result_reg_w_13[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_34 = result_reg_w_13[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_35 = result_reg_w_13[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_36 = result_reg_w_13[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_37 = result_reg_w_13[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_38 = result_reg_w_13[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_39 = result_reg_w_13[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_40 = result_reg_w_13[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_41 = result_reg_w_13[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_42 = result_reg_w_13[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_43 = result_reg_w_13[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_44 = result_reg_w_13[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_45 = result_reg_w_13[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_46 = result_reg_w_13[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_47 = result_reg_w_13[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_48 = result_reg_w_13[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_49 = result_reg_w_13[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_50 = result_reg_w_13[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_51 = result_reg_w_13[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_52 = result_reg_w_13[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_53 = result_reg_w_13[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_54 = result_reg_w_13[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_55 = result_reg_w_13[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_56 = result_reg_w_13[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_57 = result_reg_w_13[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_58 = result_reg_w_13[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_59 = result_reg_w_13[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_60 = result_reg_w_13[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_61 = result_reg_w_13[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_62 = result_reg_w_13[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_63 = result_reg_w_13[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_64 = result_reg_w_13[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_65 = result_reg_w_13[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_66 = result_reg_w_13[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_67 = result_reg_w_13[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_68 = result_reg_w_13[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_69 = result_reg_w_13[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_70 = result_reg_w_13[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_71 = result_reg_w_13[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_72 = result_reg_w_13[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_73 = result_reg_w_13[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_74 = result_reg_w_13[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_75 = result_reg_w_13[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_76 = result_reg_w_13[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_77 = result_reg_w_13[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_79 = result_reg_w_13[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_80 = result_reg_w_13[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_81 = result_reg_w_13[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_82 = result_reg_w_13[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_83 = result_reg_w_13[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_84 = result_reg_w_13[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_85 = result_reg_w_13[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_86 = result_reg_w_13[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_87 = result_reg_w_13[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_88 = result_reg_w_13[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_89 = result_reg_w_13[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_90 = result_reg_w_13[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_91 = result_reg_w_13[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_92 = result_reg_w_13[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_93 = result_reg_w_13[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_94 = result_reg_w_13[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_95 = result_reg_w_13[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_96 = result_reg_w_13[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_97 = result_reg_w_13[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_98 = result_reg_w_13[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_99 = result_reg_w_13[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_100 = result_reg_w_13[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_101 = result_reg_w_13[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_102 = result_reg_w_13[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_103 = result_reg_w_13[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_104 = result_reg_w_13[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_26_105 = result_reg_w_13[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_0 = result_reg_r_13[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_1 = result_reg_r_13[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_2 = result_reg_r_13[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_3 = result_reg_r_13[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_4 = result_reg_r_13[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_5 = result_reg_r_13[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_6 = result_reg_r_13[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_7 = result_reg_r_13[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_8 = result_reg_r_13[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_9 = result_reg_r_13[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_10 = result_reg_r_13[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_11 = result_reg_r_13[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_12 = result_reg_r_13[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_13 = result_reg_r_13[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_14 = result_reg_r_13[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_15 = result_reg_r_13[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_16 = result_reg_r_13[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_17 = result_reg_r_13[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_18 = result_reg_r_13[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_19 = result_reg_r_13[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_20 = result_reg_r_13[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_21 = result_reg_r_13[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_22 = result_reg_r_13[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_23 = result_reg_r_13[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_24 = result_reg_r_13[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_25 = result_reg_r_13[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_26 = result_reg_r_13[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_27 = result_reg_r_13[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_28 = result_reg_r_13[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_29 = result_reg_r_13[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_30 = result_reg_r_13[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_31 = result_reg_r_13[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_32 = result_reg_r_13[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_33 = result_reg_r_13[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_34 = result_reg_r_13[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_35 = result_reg_r_13[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_36 = result_reg_r_13[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_37 = result_reg_r_13[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_38 = result_reg_r_13[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_39 = result_reg_r_13[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_40 = result_reg_r_13[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_41 = result_reg_r_13[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_42 = result_reg_r_13[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_43 = result_reg_r_13[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_44 = result_reg_r_13[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_45 = result_reg_r_13[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_46 = result_reg_r_13[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_47 = result_reg_r_13[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_48 = result_reg_r_13[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_49 = result_reg_r_13[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_50 = result_reg_r_13[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_51 = result_reg_r_13[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_52 = result_reg_r_13[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_53 = result_reg_r_13[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_54 = result_reg_r_13[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_55 = result_reg_r_13[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_56 = result_reg_r_13[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_57 = result_reg_r_13[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_58 = result_reg_r_13[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_59 = result_reg_r_13[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_60 = result_reg_r_13[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_61 = result_reg_r_13[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_62 = result_reg_r_13[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_63 = result_reg_r_13[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_64 = result_reg_r_13[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_65 = result_reg_r_13[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_66 = result_reg_r_13[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_67 = result_reg_r_13[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_68 = result_reg_r_13[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_69 = result_reg_r_13[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_70 = result_reg_r_13[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_71 = result_reg_r_13[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_72 = result_reg_r_13[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_73 = result_reg_r_13[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_74 = result_reg_r_13[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_75 = result_reg_r_13[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_76 = result_reg_r_13[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_78 = result_reg_r_13[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_79 = result_reg_r_13[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_80 = result_reg_r_13[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_81 = result_reg_r_13[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_82 = result_reg_r_13[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_83 = result_reg_r_13[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_84 = result_reg_r_13[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_85 = result_reg_r_13[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_86 = result_reg_r_13[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_87 = result_reg_r_13[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_88 = result_reg_r_13[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_89 = result_reg_r_13[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_90 = result_reg_r_13[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_91 = result_reg_r_13[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_92 = result_reg_r_13[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_93 = result_reg_r_13[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_94 = result_reg_r_13[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_95 = result_reg_r_13[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_96 = result_reg_r_13[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_97 = result_reg_r_13[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_98 = result_reg_r_13[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_99 = result_reg_r_13[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_100 = result_reg_r_13[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_101 = result_reg_r_13[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_102 = result_reg_r_13[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_103 = result_reg_r_13[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_104 = result_reg_r_13[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_27_105 = result_reg_r_13[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_14_hi_hi_hi_lo = {wire_res_27_98,wire_res_27_97,wire_res_27_96,wire_res_27_95,wire_res_27_94,
    wire_res_27_93,wire_res_27_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_14_hi_hi_lo_lo = {wire_res_27_84,wire_res_27_83,wire_res_27_82,wire_res_27_81,wire_res_27_80,
    wire_res_27_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_14_hi_hi_lo = {wire_res_27_91,wire_res_27_90,wire_res_27_89,wire_res_27_88,wire_res_27_87,
    wire_res_27_86,wire_res_27_85,result_reg_w_14_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [182:0] _T_11292 = {b_aux_reg_r_13, 77'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [182:0] _GEN_1285 = {{77'd0}, a_aux_reg_r_13}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_27_77 = _GEN_1285 >= _T_11292; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_14_hi_lo_hi_lo = {wire_res_27_71,wire_res_27_70,wire_res_27_69,wire_res_27_68,wire_res_27_67,
    wire_res_27_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_14_hi_lo_lo_lo = {wire_res_27_58,wire_res_27_57,wire_res_27_56,wire_res_27_55,wire_res_27_54,
    wire_res_27_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_14_hi_lo_lo = {wire_res_27_65,wire_res_27_64,wire_res_27_63,wire_res_27_62,wire_res_27_61,
    wire_res_27_60,wire_res_27_59,result_reg_w_14_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_14_hi_lo = {wire_res_27_78,wire_res_27_77,wire_res_27_76,wire_res_27_75,wire_res_27_74,
    wire_res_27_73,wire_res_27_72,result_reg_w_14_hi_lo_hi_lo,result_reg_w_14_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_14_hi = {wire_res_27_105,wire_res_27_104,wire_res_27_103,wire_res_27_102,wire_res_27_101,
    wire_res_27_100,wire_res_27_99,result_reg_w_14_hi_hi_hi_lo,result_reg_w_14_hi_hi_lo,result_reg_w_14_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_14_lo_hi_hi_lo = {wire_res_27_45,wire_res_27_44,wire_res_27_43,wire_res_27_42,wire_res_27_41,
    wire_res_27_40,wire_res_27_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_14_lo_hi_lo_lo = {wire_res_27_31,wire_res_27_30,wire_res_27_29,wire_res_27_28,wire_res_27_27,
    wire_res_27_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_14_lo_hi_lo = {wire_res_27_38,wire_res_27_37,wire_res_27_36,wire_res_27_35,wire_res_27_34,
    wire_res_27_33,wire_res_27_32,result_reg_w_14_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_14_lo_lo_hi_lo = {wire_res_27_18,wire_res_27_17,wire_res_27_16,wire_res_27_15,wire_res_27_14,
    wire_res_27_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_14_lo_lo_lo_lo = {wire_res_27_5,wire_res_27_4,wire_res_27_3,wire_res_27_2,wire_res_27_1,
    wire_res_27_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_14_lo_lo_lo = {wire_res_27_12,wire_res_27_11,wire_res_27_10,wire_res_27_9,wire_res_27_8,
    wire_res_27_7,wire_res_27_6,result_reg_w_14_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_14_lo_lo = {wire_res_27_25,wire_res_27_24,wire_res_27_23,wire_res_27_22,wire_res_27_21,
    wire_res_27_20,wire_res_27_19,result_reg_w_14_lo_lo_hi_lo,result_reg_w_14_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_14_lo = {wire_res_27_52,wire_res_27_51,wire_res_27_50,wire_res_27_49,wire_res_27_48,
    wire_res_27_47,wire_res_27_46,result_reg_w_14_lo_hi_hi_lo,result_reg_w_14_lo_hi_lo,result_reg_w_14_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_14 = {result_reg_w_14_hi,result_reg_w_14_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_28_0 = result_reg_w_14[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_1 = result_reg_w_14[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_2 = result_reg_w_14[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_3 = result_reg_w_14[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_4 = result_reg_w_14[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_5 = result_reg_w_14[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_6 = result_reg_w_14[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_7 = result_reg_w_14[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_8 = result_reg_w_14[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_9 = result_reg_w_14[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_10 = result_reg_w_14[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_11 = result_reg_w_14[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_12 = result_reg_w_14[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_13 = result_reg_w_14[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_14 = result_reg_w_14[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_15 = result_reg_w_14[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_16 = result_reg_w_14[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_17 = result_reg_w_14[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_18 = result_reg_w_14[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_19 = result_reg_w_14[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_20 = result_reg_w_14[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_21 = result_reg_w_14[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_22 = result_reg_w_14[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_23 = result_reg_w_14[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_24 = result_reg_w_14[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_25 = result_reg_w_14[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_26 = result_reg_w_14[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_27 = result_reg_w_14[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_28 = result_reg_w_14[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_29 = result_reg_w_14[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_30 = result_reg_w_14[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_31 = result_reg_w_14[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_32 = result_reg_w_14[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_33 = result_reg_w_14[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_34 = result_reg_w_14[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_35 = result_reg_w_14[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_36 = result_reg_w_14[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_37 = result_reg_w_14[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_38 = result_reg_w_14[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_39 = result_reg_w_14[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_40 = result_reg_w_14[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_41 = result_reg_w_14[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_42 = result_reg_w_14[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_43 = result_reg_w_14[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_44 = result_reg_w_14[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_45 = result_reg_w_14[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_46 = result_reg_w_14[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_47 = result_reg_w_14[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_48 = result_reg_w_14[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_49 = result_reg_w_14[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_50 = result_reg_w_14[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_51 = result_reg_w_14[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_52 = result_reg_w_14[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_53 = result_reg_w_14[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_54 = result_reg_w_14[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_55 = result_reg_w_14[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_56 = result_reg_w_14[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_57 = result_reg_w_14[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_58 = result_reg_w_14[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_59 = result_reg_w_14[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_60 = result_reg_w_14[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_61 = result_reg_w_14[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_62 = result_reg_w_14[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_63 = result_reg_w_14[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_64 = result_reg_w_14[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_65 = result_reg_w_14[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_66 = result_reg_w_14[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_67 = result_reg_w_14[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_68 = result_reg_w_14[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_69 = result_reg_w_14[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_70 = result_reg_w_14[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_71 = result_reg_w_14[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_72 = result_reg_w_14[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_73 = result_reg_w_14[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_74 = result_reg_w_14[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_75 = result_reg_w_14[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_77 = result_reg_w_14[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_78 = result_reg_w_14[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_79 = result_reg_w_14[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_80 = result_reg_w_14[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_81 = result_reg_w_14[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_82 = result_reg_w_14[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_83 = result_reg_w_14[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_84 = result_reg_w_14[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_85 = result_reg_w_14[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_86 = result_reg_w_14[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_87 = result_reg_w_14[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_88 = result_reg_w_14[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_89 = result_reg_w_14[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_90 = result_reg_w_14[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_91 = result_reg_w_14[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_92 = result_reg_w_14[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_93 = result_reg_w_14[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_94 = result_reg_w_14[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_95 = result_reg_w_14[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_96 = result_reg_w_14[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_97 = result_reg_w_14[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_98 = result_reg_w_14[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_99 = result_reg_w_14[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_100 = result_reg_w_14[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_101 = result_reg_w_14[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_102 = result_reg_w_14[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_103 = result_reg_w_14[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_104 = result_reg_w_14[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_28_105 = result_reg_w_14[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_0 = result_reg_r_14[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_1 = result_reg_r_14[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_2 = result_reg_r_14[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_3 = result_reg_r_14[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_4 = result_reg_r_14[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_5 = result_reg_r_14[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_6 = result_reg_r_14[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_7 = result_reg_r_14[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_8 = result_reg_r_14[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_9 = result_reg_r_14[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_10 = result_reg_r_14[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_11 = result_reg_r_14[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_12 = result_reg_r_14[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_13 = result_reg_r_14[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_14 = result_reg_r_14[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_15 = result_reg_r_14[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_16 = result_reg_r_14[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_17 = result_reg_r_14[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_18 = result_reg_r_14[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_19 = result_reg_r_14[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_20 = result_reg_r_14[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_21 = result_reg_r_14[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_22 = result_reg_r_14[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_23 = result_reg_r_14[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_24 = result_reg_r_14[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_25 = result_reg_r_14[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_26 = result_reg_r_14[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_27 = result_reg_r_14[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_28 = result_reg_r_14[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_29 = result_reg_r_14[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_30 = result_reg_r_14[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_31 = result_reg_r_14[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_32 = result_reg_r_14[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_33 = result_reg_r_14[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_34 = result_reg_r_14[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_35 = result_reg_r_14[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_36 = result_reg_r_14[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_37 = result_reg_r_14[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_38 = result_reg_r_14[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_39 = result_reg_r_14[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_40 = result_reg_r_14[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_41 = result_reg_r_14[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_42 = result_reg_r_14[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_43 = result_reg_r_14[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_44 = result_reg_r_14[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_45 = result_reg_r_14[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_46 = result_reg_r_14[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_47 = result_reg_r_14[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_48 = result_reg_r_14[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_49 = result_reg_r_14[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_50 = result_reg_r_14[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_51 = result_reg_r_14[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_52 = result_reg_r_14[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_53 = result_reg_r_14[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_54 = result_reg_r_14[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_55 = result_reg_r_14[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_56 = result_reg_r_14[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_57 = result_reg_r_14[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_58 = result_reg_r_14[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_59 = result_reg_r_14[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_60 = result_reg_r_14[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_61 = result_reg_r_14[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_62 = result_reg_r_14[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_63 = result_reg_r_14[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_64 = result_reg_r_14[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_65 = result_reg_r_14[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_66 = result_reg_r_14[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_67 = result_reg_r_14[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_68 = result_reg_r_14[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_69 = result_reg_r_14[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_70 = result_reg_r_14[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_71 = result_reg_r_14[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_72 = result_reg_r_14[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_73 = result_reg_r_14[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_74 = result_reg_r_14[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_76 = result_reg_r_14[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_77 = result_reg_r_14[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_78 = result_reg_r_14[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_79 = result_reg_r_14[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_80 = result_reg_r_14[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_81 = result_reg_r_14[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_82 = result_reg_r_14[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_83 = result_reg_r_14[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_84 = result_reg_r_14[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_85 = result_reg_r_14[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_86 = result_reg_r_14[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_87 = result_reg_r_14[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_88 = result_reg_r_14[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_89 = result_reg_r_14[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_90 = result_reg_r_14[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_91 = result_reg_r_14[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_92 = result_reg_r_14[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_93 = result_reg_r_14[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_94 = result_reg_r_14[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_95 = result_reg_r_14[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_96 = result_reg_r_14[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_97 = result_reg_r_14[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_98 = result_reg_r_14[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_99 = result_reg_r_14[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_100 = result_reg_r_14[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_101 = result_reg_r_14[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_102 = result_reg_r_14[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_103 = result_reg_r_14[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_104 = result_reg_r_14[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_29_105 = result_reg_r_14[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_15_hi_hi_hi_lo = {wire_res_29_98,wire_res_29_97,wire_res_29_96,wire_res_29_95,wire_res_29_94,
    wire_res_29_93,wire_res_29_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_15_hi_hi_lo_lo = {wire_res_29_84,wire_res_29_83,wire_res_29_82,wire_res_29_81,wire_res_29_80,
    wire_res_29_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_15_hi_hi_lo = {wire_res_29_91,wire_res_29_90,wire_res_29_89,wire_res_29_88,wire_res_29_87,
    wire_res_29_86,wire_res_29_85,result_reg_w_15_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [180:0] _T_11296 = {b_aux_reg_r_14, 75'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [180:0] _GEN_1286 = {{75'd0}, a_aux_reg_r_14}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_29_75 = _GEN_1286 >= _T_11296; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_15_hi_lo_hi_lo = {wire_res_29_71,wire_res_29_70,wire_res_29_69,wire_res_29_68,wire_res_29_67,
    wire_res_29_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_15_hi_lo_lo_lo = {wire_res_29_58,wire_res_29_57,wire_res_29_56,wire_res_29_55,wire_res_29_54,
    wire_res_29_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_15_hi_lo_lo = {wire_res_29_65,wire_res_29_64,wire_res_29_63,wire_res_29_62,wire_res_29_61,
    wire_res_29_60,wire_res_29_59,result_reg_w_15_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_15_hi_lo = {wire_res_29_78,wire_res_29_77,wire_res_29_76,wire_res_29_75,wire_res_29_74,
    wire_res_29_73,wire_res_29_72,result_reg_w_15_hi_lo_hi_lo,result_reg_w_15_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_15_hi = {wire_res_29_105,wire_res_29_104,wire_res_29_103,wire_res_29_102,wire_res_29_101,
    wire_res_29_100,wire_res_29_99,result_reg_w_15_hi_hi_hi_lo,result_reg_w_15_hi_hi_lo,result_reg_w_15_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_15_lo_hi_hi_lo = {wire_res_29_45,wire_res_29_44,wire_res_29_43,wire_res_29_42,wire_res_29_41,
    wire_res_29_40,wire_res_29_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_15_lo_hi_lo_lo = {wire_res_29_31,wire_res_29_30,wire_res_29_29,wire_res_29_28,wire_res_29_27,
    wire_res_29_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_15_lo_hi_lo = {wire_res_29_38,wire_res_29_37,wire_res_29_36,wire_res_29_35,wire_res_29_34,
    wire_res_29_33,wire_res_29_32,result_reg_w_15_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_15_lo_lo_hi_lo = {wire_res_29_18,wire_res_29_17,wire_res_29_16,wire_res_29_15,wire_res_29_14,
    wire_res_29_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_15_lo_lo_lo_lo = {wire_res_29_5,wire_res_29_4,wire_res_29_3,wire_res_29_2,wire_res_29_1,
    wire_res_29_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_15_lo_lo_lo = {wire_res_29_12,wire_res_29_11,wire_res_29_10,wire_res_29_9,wire_res_29_8,
    wire_res_29_7,wire_res_29_6,result_reg_w_15_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_15_lo_lo = {wire_res_29_25,wire_res_29_24,wire_res_29_23,wire_res_29_22,wire_res_29_21,
    wire_res_29_20,wire_res_29_19,result_reg_w_15_lo_lo_hi_lo,result_reg_w_15_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_15_lo = {wire_res_29_52,wire_res_29_51,wire_res_29_50,wire_res_29_49,wire_res_29_48,
    wire_res_29_47,wire_res_29_46,result_reg_w_15_lo_hi_hi_lo,result_reg_w_15_lo_hi_lo,result_reg_w_15_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_15 = {result_reg_w_15_hi,result_reg_w_15_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_30_0 = result_reg_w_15[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_1 = result_reg_w_15[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_2 = result_reg_w_15[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_3 = result_reg_w_15[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_4 = result_reg_w_15[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_5 = result_reg_w_15[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_6 = result_reg_w_15[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_7 = result_reg_w_15[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_8 = result_reg_w_15[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_9 = result_reg_w_15[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_10 = result_reg_w_15[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_11 = result_reg_w_15[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_12 = result_reg_w_15[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_13 = result_reg_w_15[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_14 = result_reg_w_15[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_15 = result_reg_w_15[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_16 = result_reg_w_15[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_17 = result_reg_w_15[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_18 = result_reg_w_15[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_19 = result_reg_w_15[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_20 = result_reg_w_15[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_21 = result_reg_w_15[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_22 = result_reg_w_15[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_23 = result_reg_w_15[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_24 = result_reg_w_15[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_25 = result_reg_w_15[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_26 = result_reg_w_15[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_27 = result_reg_w_15[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_28 = result_reg_w_15[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_29 = result_reg_w_15[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_30 = result_reg_w_15[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_31 = result_reg_w_15[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_32 = result_reg_w_15[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_33 = result_reg_w_15[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_34 = result_reg_w_15[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_35 = result_reg_w_15[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_36 = result_reg_w_15[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_37 = result_reg_w_15[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_38 = result_reg_w_15[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_39 = result_reg_w_15[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_40 = result_reg_w_15[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_41 = result_reg_w_15[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_42 = result_reg_w_15[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_43 = result_reg_w_15[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_44 = result_reg_w_15[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_45 = result_reg_w_15[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_46 = result_reg_w_15[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_47 = result_reg_w_15[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_48 = result_reg_w_15[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_49 = result_reg_w_15[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_50 = result_reg_w_15[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_51 = result_reg_w_15[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_52 = result_reg_w_15[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_53 = result_reg_w_15[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_54 = result_reg_w_15[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_55 = result_reg_w_15[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_56 = result_reg_w_15[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_57 = result_reg_w_15[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_58 = result_reg_w_15[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_59 = result_reg_w_15[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_60 = result_reg_w_15[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_61 = result_reg_w_15[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_62 = result_reg_w_15[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_63 = result_reg_w_15[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_64 = result_reg_w_15[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_65 = result_reg_w_15[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_66 = result_reg_w_15[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_67 = result_reg_w_15[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_68 = result_reg_w_15[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_69 = result_reg_w_15[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_70 = result_reg_w_15[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_71 = result_reg_w_15[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_72 = result_reg_w_15[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_73 = result_reg_w_15[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_75 = result_reg_w_15[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_76 = result_reg_w_15[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_77 = result_reg_w_15[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_78 = result_reg_w_15[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_79 = result_reg_w_15[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_80 = result_reg_w_15[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_81 = result_reg_w_15[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_82 = result_reg_w_15[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_83 = result_reg_w_15[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_84 = result_reg_w_15[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_85 = result_reg_w_15[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_86 = result_reg_w_15[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_87 = result_reg_w_15[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_88 = result_reg_w_15[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_89 = result_reg_w_15[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_90 = result_reg_w_15[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_91 = result_reg_w_15[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_92 = result_reg_w_15[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_93 = result_reg_w_15[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_94 = result_reg_w_15[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_95 = result_reg_w_15[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_96 = result_reg_w_15[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_97 = result_reg_w_15[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_98 = result_reg_w_15[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_99 = result_reg_w_15[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_100 = result_reg_w_15[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_101 = result_reg_w_15[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_102 = result_reg_w_15[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_103 = result_reg_w_15[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_104 = result_reg_w_15[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_30_105 = result_reg_w_15[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_0 = result_reg_r_15[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_1 = result_reg_r_15[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_2 = result_reg_r_15[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_3 = result_reg_r_15[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_4 = result_reg_r_15[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_5 = result_reg_r_15[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_6 = result_reg_r_15[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_7 = result_reg_r_15[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_8 = result_reg_r_15[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_9 = result_reg_r_15[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_10 = result_reg_r_15[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_11 = result_reg_r_15[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_12 = result_reg_r_15[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_13 = result_reg_r_15[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_14 = result_reg_r_15[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_15 = result_reg_r_15[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_16 = result_reg_r_15[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_17 = result_reg_r_15[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_18 = result_reg_r_15[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_19 = result_reg_r_15[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_20 = result_reg_r_15[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_21 = result_reg_r_15[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_22 = result_reg_r_15[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_23 = result_reg_r_15[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_24 = result_reg_r_15[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_25 = result_reg_r_15[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_26 = result_reg_r_15[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_27 = result_reg_r_15[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_28 = result_reg_r_15[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_29 = result_reg_r_15[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_30 = result_reg_r_15[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_31 = result_reg_r_15[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_32 = result_reg_r_15[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_33 = result_reg_r_15[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_34 = result_reg_r_15[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_35 = result_reg_r_15[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_36 = result_reg_r_15[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_37 = result_reg_r_15[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_38 = result_reg_r_15[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_39 = result_reg_r_15[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_40 = result_reg_r_15[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_41 = result_reg_r_15[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_42 = result_reg_r_15[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_43 = result_reg_r_15[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_44 = result_reg_r_15[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_45 = result_reg_r_15[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_46 = result_reg_r_15[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_47 = result_reg_r_15[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_48 = result_reg_r_15[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_49 = result_reg_r_15[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_50 = result_reg_r_15[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_51 = result_reg_r_15[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_52 = result_reg_r_15[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_53 = result_reg_r_15[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_54 = result_reg_r_15[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_55 = result_reg_r_15[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_56 = result_reg_r_15[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_57 = result_reg_r_15[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_58 = result_reg_r_15[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_59 = result_reg_r_15[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_60 = result_reg_r_15[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_61 = result_reg_r_15[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_62 = result_reg_r_15[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_63 = result_reg_r_15[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_64 = result_reg_r_15[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_65 = result_reg_r_15[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_66 = result_reg_r_15[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_67 = result_reg_r_15[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_68 = result_reg_r_15[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_69 = result_reg_r_15[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_70 = result_reg_r_15[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_71 = result_reg_r_15[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_72 = result_reg_r_15[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_74 = result_reg_r_15[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_75 = result_reg_r_15[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_76 = result_reg_r_15[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_77 = result_reg_r_15[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_78 = result_reg_r_15[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_79 = result_reg_r_15[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_80 = result_reg_r_15[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_81 = result_reg_r_15[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_82 = result_reg_r_15[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_83 = result_reg_r_15[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_84 = result_reg_r_15[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_85 = result_reg_r_15[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_86 = result_reg_r_15[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_87 = result_reg_r_15[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_88 = result_reg_r_15[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_89 = result_reg_r_15[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_90 = result_reg_r_15[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_91 = result_reg_r_15[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_92 = result_reg_r_15[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_93 = result_reg_r_15[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_94 = result_reg_r_15[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_95 = result_reg_r_15[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_96 = result_reg_r_15[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_97 = result_reg_r_15[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_98 = result_reg_r_15[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_99 = result_reg_r_15[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_100 = result_reg_r_15[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_101 = result_reg_r_15[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_102 = result_reg_r_15[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_103 = result_reg_r_15[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_104 = result_reg_r_15[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_31_105 = result_reg_r_15[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_16_hi_hi_hi_lo = {wire_res_31_98,wire_res_31_97,wire_res_31_96,wire_res_31_95,wire_res_31_94,
    wire_res_31_93,wire_res_31_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_16_hi_hi_lo_lo = {wire_res_31_84,wire_res_31_83,wire_res_31_82,wire_res_31_81,wire_res_31_80,
    wire_res_31_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_16_hi_hi_lo = {wire_res_31_91,wire_res_31_90,wire_res_31_89,wire_res_31_88,wire_res_31_87,
    wire_res_31_86,wire_res_31_85,result_reg_w_16_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [178:0] _T_11300 = {b_aux_reg_r_15, 73'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [178:0] _GEN_1287 = {{73'd0}, a_aux_reg_r_15}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_31_73 = _GEN_1287 >= _T_11300; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_16_hi_lo_hi_lo = {wire_res_31_71,wire_res_31_70,wire_res_31_69,wire_res_31_68,wire_res_31_67,
    wire_res_31_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_16_hi_lo_lo_lo = {wire_res_31_58,wire_res_31_57,wire_res_31_56,wire_res_31_55,wire_res_31_54,
    wire_res_31_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_16_hi_lo_lo = {wire_res_31_65,wire_res_31_64,wire_res_31_63,wire_res_31_62,wire_res_31_61,
    wire_res_31_60,wire_res_31_59,result_reg_w_16_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_16_hi_lo = {wire_res_31_78,wire_res_31_77,wire_res_31_76,wire_res_31_75,wire_res_31_74,
    wire_res_31_73,wire_res_31_72,result_reg_w_16_hi_lo_hi_lo,result_reg_w_16_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_16_hi = {wire_res_31_105,wire_res_31_104,wire_res_31_103,wire_res_31_102,wire_res_31_101,
    wire_res_31_100,wire_res_31_99,result_reg_w_16_hi_hi_hi_lo,result_reg_w_16_hi_hi_lo,result_reg_w_16_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_16_lo_hi_hi_lo = {wire_res_31_45,wire_res_31_44,wire_res_31_43,wire_res_31_42,wire_res_31_41,
    wire_res_31_40,wire_res_31_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_16_lo_hi_lo_lo = {wire_res_31_31,wire_res_31_30,wire_res_31_29,wire_res_31_28,wire_res_31_27,
    wire_res_31_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_16_lo_hi_lo = {wire_res_31_38,wire_res_31_37,wire_res_31_36,wire_res_31_35,wire_res_31_34,
    wire_res_31_33,wire_res_31_32,result_reg_w_16_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_16_lo_lo_hi_lo = {wire_res_31_18,wire_res_31_17,wire_res_31_16,wire_res_31_15,wire_res_31_14,
    wire_res_31_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_16_lo_lo_lo_lo = {wire_res_31_5,wire_res_31_4,wire_res_31_3,wire_res_31_2,wire_res_31_1,
    wire_res_31_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_16_lo_lo_lo = {wire_res_31_12,wire_res_31_11,wire_res_31_10,wire_res_31_9,wire_res_31_8,
    wire_res_31_7,wire_res_31_6,result_reg_w_16_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_16_lo_lo = {wire_res_31_25,wire_res_31_24,wire_res_31_23,wire_res_31_22,wire_res_31_21,
    wire_res_31_20,wire_res_31_19,result_reg_w_16_lo_lo_hi_lo,result_reg_w_16_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_16_lo = {wire_res_31_52,wire_res_31_51,wire_res_31_50,wire_res_31_49,wire_res_31_48,
    wire_res_31_47,wire_res_31_46,result_reg_w_16_lo_hi_hi_lo,result_reg_w_16_lo_hi_lo,result_reg_w_16_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_16 = {result_reg_w_16_hi,result_reg_w_16_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_32_0 = result_reg_w_16[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_1 = result_reg_w_16[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_2 = result_reg_w_16[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_3 = result_reg_w_16[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_4 = result_reg_w_16[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_5 = result_reg_w_16[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_6 = result_reg_w_16[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_7 = result_reg_w_16[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_8 = result_reg_w_16[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_9 = result_reg_w_16[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_10 = result_reg_w_16[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_11 = result_reg_w_16[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_12 = result_reg_w_16[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_13 = result_reg_w_16[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_14 = result_reg_w_16[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_15 = result_reg_w_16[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_16 = result_reg_w_16[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_17 = result_reg_w_16[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_18 = result_reg_w_16[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_19 = result_reg_w_16[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_20 = result_reg_w_16[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_21 = result_reg_w_16[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_22 = result_reg_w_16[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_23 = result_reg_w_16[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_24 = result_reg_w_16[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_25 = result_reg_w_16[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_26 = result_reg_w_16[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_27 = result_reg_w_16[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_28 = result_reg_w_16[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_29 = result_reg_w_16[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_30 = result_reg_w_16[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_31 = result_reg_w_16[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_32 = result_reg_w_16[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_33 = result_reg_w_16[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_34 = result_reg_w_16[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_35 = result_reg_w_16[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_36 = result_reg_w_16[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_37 = result_reg_w_16[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_38 = result_reg_w_16[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_39 = result_reg_w_16[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_40 = result_reg_w_16[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_41 = result_reg_w_16[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_42 = result_reg_w_16[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_43 = result_reg_w_16[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_44 = result_reg_w_16[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_45 = result_reg_w_16[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_46 = result_reg_w_16[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_47 = result_reg_w_16[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_48 = result_reg_w_16[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_49 = result_reg_w_16[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_50 = result_reg_w_16[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_51 = result_reg_w_16[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_52 = result_reg_w_16[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_53 = result_reg_w_16[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_54 = result_reg_w_16[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_55 = result_reg_w_16[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_56 = result_reg_w_16[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_57 = result_reg_w_16[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_58 = result_reg_w_16[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_59 = result_reg_w_16[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_60 = result_reg_w_16[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_61 = result_reg_w_16[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_62 = result_reg_w_16[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_63 = result_reg_w_16[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_64 = result_reg_w_16[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_65 = result_reg_w_16[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_66 = result_reg_w_16[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_67 = result_reg_w_16[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_68 = result_reg_w_16[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_69 = result_reg_w_16[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_70 = result_reg_w_16[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_71 = result_reg_w_16[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_73 = result_reg_w_16[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_74 = result_reg_w_16[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_75 = result_reg_w_16[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_76 = result_reg_w_16[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_77 = result_reg_w_16[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_78 = result_reg_w_16[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_79 = result_reg_w_16[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_80 = result_reg_w_16[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_81 = result_reg_w_16[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_82 = result_reg_w_16[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_83 = result_reg_w_16[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_84 = result_reg_w_16[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_85 = result_reg_w_16[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_86 = result_reg_w_16[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_87 = result_reg_w_16[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_88 = result_reg_w_16[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_89 = result_reg_w_16[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_90 = result_reg_w_16[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_91 = result_reg_w_16[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_92 = result_reg_w_16[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_93 = result_reg_w_16[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_94 = result_reg_w_16[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_95 = result_reg_w_16[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_96 = result_reg_w_16[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_97 = result_reg_w_16[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_98 = result_reg_w_16[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_99 = result_reg_w_16[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_100 = result_reg_w_16[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_101 = result_reg_w_16[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_102 = result_reg_w_16[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_103 = result_reg_w_16[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_104 = result_reg_w_16[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_32_105 = result_reg_w_16[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_0 = result_reg_r_16[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_1 = result_reg_r_16[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_2 = result_reg_r_16[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_3 = result_reg_r_16[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_4 = result_reg_r_16[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_5 = result_reg_r_16[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_6 = result_reg_r_16[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_7 = result_reg_r_16[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_8 = result_reg_r_16[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_9 = result_reg_r_16[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_10 = result_reg_r_16[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_11 = result_reg_r_16[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_12 = result_reg_r_16[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_13 = result_reg_r_16[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_14 = result_reg_r_16[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_15 = result_reg_r_16[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_16 = result_reg_r_16[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_17 = result_reg_r_16[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_18 = result_reg_r_16[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_19 = result_reg_r_16[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_20 = result_reg_r_16[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_21 = result_reg_r_16[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_22 = result_reg_r_16[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_23 = result_reg_r_16[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_24 = result_reg_r_16[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_25 = result_reg_r_16[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_26 = result_reg_r_16[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_27 = result_reg_r_16[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_28 = result_reg_r_16[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_29 = result_reg_r_16[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_30 = result_reg_r_16[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_31 = result_reg_r_16[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_32 = result_reg_r_16[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_33 = result_reg_r_16[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_34 = result_reg_r_16[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_35 = result_reg_r_16[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_36 = result_reg_r_16[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_37 = result_reg_r_16[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_38 = result_reg_r_16[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_39 = result_reg_r_16[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_40 = result_reg_r_16[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_41 = result_reg_r_16[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_42 = result_reg_r_16[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_43 = result_reg_r_16[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_44 = result_reg_r_16[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_45 = result_reg_r_16[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_46 = result_reg_r_16[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_47 = result_reg_r_16[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_48 = result_reg_r_16[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_49 = result_reg_r_16[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_50 = result_reg_r_16[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_51 = result_reg_r_16[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_52 = result_reg_r_16[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_53 = result_reg_r_16[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_54 = result_reg_r_16[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_55 = result_reg_r_16[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_56 = result_reg_r_16[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_57 = result_reg_r_16[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_58 = result_reg_r_16[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_59 = result_reg_r_16[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_60 = result_reg_r_16[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_61 = result_reg_r_16[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_62 = result_reg_r_16[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_63 = result_reg_r_16[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_64 = result_reg_r_16[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_65 = result_reg_r_16[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_66 = result_reg_r_16[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_67 = result_reg_r_16[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_68 = result_reg_r_16[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_69 = result_reg_r_16[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_70 = result_reg_r_16[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_72 = result_reg_r_16[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_73 = result_reg_r_16[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_74 = result_reg_r_16[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_75 = result_reg_r_16[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_76 = result_reg_r_16[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_77 = result_reg_r_16[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_78 = result_reg_r_16[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_79 = result_reg_r_16[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_80 = result_reg_r_16[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_81 = result_reg_r_16[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_82 = result_reg_r_16[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_83 = result_reg_r_16[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_84 = result_reg_r_16[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_85 = result_reg_r_16[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_86 = result_reg_r_16[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_87 = result_reg_r_16[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_88 = result_reg_r_16[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_89 = result_reg_r_16[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_90 = result_reg_r_16[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_91 = result_reg_r_16[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_92 = result_reg_r_16[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_93 = result_reg_r_16[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_94 = result_reg_r_16[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_95 = result_reg_r_16[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_96 = result_reg_r_16[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_97 = result_reg_r_16[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_98 = result_reg_r_16[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_99 = result_reg_r_16[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_100 = result_reg_r_16[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_101 = result_reg_r_16[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_102 = result_reg_r_16[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_103 = result_reg_r_16[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_104 = result_reg_r_16[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_33_105 = result_reg_r_16[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_17_hi_hi_hi_lo = {wire_res_33_98,wire_res_33_97,wire_res_33_96,wire_res_33_95,wire_res_33_94,
    wire_res_33_93,wire_res_33_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_17_hi_hi_lo_lo = {wire_res_33_84,wire_res_33_83,wire_res_33_82,wire_res_33_81,wire_res_33_80,
    wire_res_33_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_17_hi_hi_lo = {wire_res_33_91,wire_res_33_90,wire_res_33_89,wire_res_33_88,wire_res_33_87,
    wire_res_33_86,wire_res_33_85,result_reg_w_17_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [176:0] _T_11304 = {b_aux_reg_r_16, 71'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [176:0] _GEN_1288 = {{71'd0}, a_aux_reg_r_16}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_33_71 = _GEN_1288 >= _T_11304; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_17_hi_lo_hi_lo = {wire_res_33_71,wire_res_33_70,wire_res_33_69,wire_res_33_68,wire_res_33_67,
    wire_res_33_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_17_hi_lo_lo_lo = {wire_res_33_58,wire_res_33_57,wire_res_33_56,wire_res_33_55,wire_res_33_54,
    wire_res_33_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_17_hi_lo_lo = {wire_res_33_65,wire_res_33_64,wire_res_33_63,wire_res_33_62,wire_res_33_61,
    wire_res_33_60,wire_res_33_59,result_reg_w_17_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_17_hi_lo = {wire_res_33_78,wire_res_33_77,wire_res_33_76,wire_res_33_75,wire_res_33_74,
    wire_res_33_73,wire_res_33_72,result_reg_w_17_hi_lo_hi_lo,result_reg_w_17_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_17_hi = {wire_res_33_105,wire_res_33_104,wire_res_33_103,wire_res_33_102,wire_res_33_101,
    wire_res_33_100,wire_res_33_99,result_reg_w_17_hi_hi_hi_lo,result_reg_w_17_hi_hi_lo,result_reg_w_17_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_17_lo_hi_hi_lo = {wire_res_33_45,wire_res_33_44,wire_res_33_43,wire_res_33_42,wire_res_33_41,
    wire_res_33_40,wire_res_33_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_17_lo_hi_lo_lo = {wire_res_33_31,wire_res_33_30,wire_res_33_29,wire_res_33_28,wire_res_33_27,
    wire_res_33_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_17_lo_hi_lo = {wire_res_33_38,wire_res_33_37,wire_res_33_36,wire_res_33_35,wire_res_33_34,
    wire_res_33_33,wire_res_33_32,result_reg_w_17_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_17_lo_lo_hi_lo = {wire_res_33_18,wire_res_33_17,wire_res_33_16,wire_res_33_15,wire_res_33_14,
    wire_res_33_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_17_lo_lo_lo_lo = {wire_res_33_5,wire_res_33_4,wire_res_33_3,wire_res_33_2,wire_res_33_1,
    wire_res_33_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_17_lo_lo_lo = {wire_res_33_12,wire_res_33_11,wire_res_33_10,wire_res_33_9,wire_res_33_8,
    wire_res_33_7,wire_res_33_6,result_reg_w_17_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_17_lo_lo = {wire_res_33_25,wire_res_33_24,wire_res_33_23,wire_res_33_22,wire_res_33_21,
    wire_res_33_20,wire_res_33_19,result_reg_w_17_lo_lo_hi_lo,result_reg_w_17_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_17_lo = {wire_res_33_52,wire_res_33_51,wire_res_33_50,wire_res_33_49,wire_res_33_48,
    wire_res_33_47,wire_res_33_46,result_reg_w_17_lo_hi_hi_lo,result_reg_w_17_lo_hi_lo,result_reg_w_17_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_17 = {result_reg_w_17_hi,result_reg_w_17_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_34_0 = result_reg_w_17[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_1 = result_reg_w_17[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_2 = result_reg_w_17[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_3 = result_reg_w_17[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_4 = result_reg_w_17[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_5 = result_reg_w_17[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_6 = result_reg_w_17[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_7 = result_reg_w_17[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_8 = result_reg_w_17[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_9 = result_reg_w_17[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_10 = result_reg_w_17[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_11 = result_reg_w_17[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_12 = result_reg_w_17[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_13 = result_reg_w_17[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_14 = result_reg_w_17[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_15 = result_reg_w_17[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_16 = result_reg_w_17[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_17 = result_reg_w_17[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_18 = result_reg_w_17[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_19 = result_reg_w_17[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_20 = result_reg_w_17[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_21 = result_reg_w_17[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_22 = result_reg_w_17[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_23 = result_reg_w_17[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_24 = result_reg_w_17[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_25 = result_reg_w_17[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_26 = result_reg_w_17[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_27 = result_reg_w_17[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_28 = result_reg_w_17[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_29 = result_reg_w_17[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_30 = result_reg_w_17[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_31 = result_reg_w_17[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_32 = result_reg_w_17[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_33 = result_reg_w_17[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_34 = result_reg_w_17[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_35 = result_reg_w_17[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_36 = result_reg_w_17[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_37 = result_reg_w_17[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_38 = result_reg_w_17[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_39 = result_reg_w_17[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_40 = result_reg_w_17[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_41 = result_reg_w_17[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_42 = result_reg_w_17[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_43 = result_reg_w_17[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_44 = result_reg_w_17[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_45 = result_reg_w_17[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_46 = result_reg_w_17[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_47 = result_reg_w_17[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_48 = result_reg_w_17[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_49 = result_reg_w_17[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_50 = result_reg_w_17[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_51 = result_reg_w_17[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_52 = result_reg_w_17[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_53 = result_reg_w_17[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_54 = result_reg_w_17[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_55 = result_reg_w_17[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_56 = result_reg_w_17[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_57 = result_reg_w_17[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_58 = result_reg_w_17[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_59 = result_reg_w_17[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_60 = result_reg_w_17[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_61 = result_reg_w_17[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_62 = result_reg_w_17[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_63 = result_reg_w_17[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_64 = result_reg_w_17[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_65 = result_reg_w_17[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_66 = result_reg_w_17[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_67 = result_reg_w_17[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_68 = result_reg_w_17[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_69 = result_reg_w_17[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_71 = result_reg_w_17[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_72 = result_reg_w_17[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_73 = result_reg_w_17[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_74 = result_reg_w_17[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_75 = result_reg_w_17[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_76 = result_reg_w_17[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_77 = result_reg_w_17[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_78 = result_reg_w_17[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_79 = result_reg_w_17[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_80 = result_reg_w_17[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_81 = result_reg_w_17[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_82 = result_reg_w_17[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_83 = result_reg_w_17[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_84 = result_reg_w_17[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_85 = result_reg_w_17[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_86 = result_reg_w_17[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_87 = result_reg_w_17[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_88 = result_reg_w_17[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_89 = result_reg_w_17[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_90 = result_reg_w_17[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_91 = result_reg_w_17[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_92 = result_reg_w_17[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_93 = result_reg_w_17[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_94 = result_reg_w_17[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_95 = result_reg_w_17[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_96 = result_reg_w_17[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_97 = result_reg_w_17[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_98 = result_reg_w_17[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_99 = result_reg_w_17[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_100 = result_reg_w_17[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_101 = result_reg_w_17[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_102 = result_reg_w_17[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_103 = result_reg_w_17[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_104 = result_reg_w_17[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_34_105 = result_reg_w_17[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_0 = result_reg_r_17[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_1 = result_reg_r_17[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_2 = result_reg_r_17[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_3 = result_reg_r_17[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_4 = result_reg_r_17[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_5 = result_reg_r_17[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_6 = result_reg_r_17[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_7 = result_reg_r_17[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_8 = result_reg_r_17[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_9 = result_reg_r_17[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_10 = result_reg_r_17[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_11 = result_reg_r_17[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_12 = result_reg_r_17[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_13 = result_reg_r_17[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_14 = result_reg_r_17[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_15 = result_reg_r_17[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_16 = result_reg_r_17[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_17 = result_reg_r_17[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_18 = result_reg_r_17[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_19 = result_reg_r_17[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_20 = result_reg_r_17[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_21 = result_reg_r_17[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_22 = result_reg_r_17[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_23 = result_reg_r_17[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_24 = result_reg_r_17[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_25 = result_reg_r_17[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_26 = result_reg_r_17[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_27 = result_reg_r_17[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_28 = result_reg_r_17[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_29 = result_reg_r_17[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_30 = result_reg_r_17[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_31 = result_reg_r_17[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_32 = result_reg_r_17[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_33 = result_reg_r_17[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_34 = result_reg_r_17[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_35 = result_reg_r_17[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_36 = result_reg_r_17[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_37 = result_reg_r_17[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_38 = result_reg_r_17[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_39 = result_reg_r_17[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_40 = result_reg_r_17[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_41 = result_reg_r_17[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_42 = result_reg_r_17[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_43 = result_reg_r_17[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_44 = result_reg_r_17[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_45 = result_reg_r_17[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_46 = result_reg_r_17[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_47 = result_reg_r_17[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_48 = result_reg_r_17[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_49 = result_reg_r_17[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_50 = result_reg_r_17[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_51 = result_reg_r_17[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_52 = result_reg_r_17[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_53 = result_reg_r_17[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_54 = result_reg_r_17[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_55 = result_reg_r_17[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_56 = result_reg_r_17[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_57 = result_reg_r_17[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_58 = result_reg_r_17[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_59 = result_reg_r_17[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_60 = result_reg_r_17[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_61 = result_reg_r_17[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_62 = result_reg_r_17[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_63 = result_reg_r_17[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_64 = result_reg_r_17[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_65 = result_reg_r_17[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_66 = result_reg_r_17[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_67 = result_reg_r_17[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_68 = result_reg_r_17[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_70 = result_reg_r_17[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_71 = result_reg_r_17[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_72 = result_reg_r_17[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_73 = result_reg_r_17[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_74 = result_reg_r_17[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_75 = result_reg_r_17[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_76 = result_reg_r_17[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_77 = result_reg_r_17[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_78 = result_reg_r_17[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_79 = result_reg_r_17[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_80 = result_reg_r_17[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_81 = result_reg_r_17[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_82 = result_reg_r_17[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_83 = result_reg_r_17[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_84 = result_reg_r_17[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_85 = result_reg_r_17[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_86 = result_reg_r_17[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_87 = result_reg_r_17[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_88 = result_reg_r_17[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_89 = result_reg_r_17[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_90 = result_reg_r_17[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_91 = result_reg_r_17[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_92 = result_reg_r_17[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_93 = result_reg_r_17[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_94 = result_reg_r_17[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_95 = result_reg_r_17[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_96 = result_reg_r_17[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_97 = result_reg_r_17[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_98 = result_reg_r_17[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_99 = result_reg_r_17[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_100 = result_reg_r_17[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_101 = result_reg_r_17[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_102 = result_reg_r_17[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_103 = result_reg_r_17[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_104 = result_reg_r_17[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_35_105 = result_reg_r_17[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_18_hi_hi_hi_lo = {wire_res_35_98,wire_res_35_97,wire_res_35_96,wire_res_35_95,wire_res_35_94,
    wire_res_35_93,wire_res_35_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_18_hi_hi_lo_lo = {wire_res_35_84,wire_res_35_83,wire_res_35_82,wire_res_35_81,wire_res_35_80,
    wire_res_35_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_18_hi_hi_lo = {wire_res_35_91,wire_res_35_90,wire_res_35_89,wire_res_35_88,wire_res_35_87,
    wire_res_35_86,wire_res_35_85,result_reg_w_18_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [174:0] _T_11308 = {b_aux_reg_r_17, 69'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [174:0] _GEN_1289 = {{69'd0}, a_aux_reg_r_17}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_35_69 = _GEN_1289 >= _T_11308; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_18_hi_lo_hi_lo = {wire_res_35_71,wire_res_35_70,wire_res_35_69,wire_res_35_68,wire_res_35_67,
    wire_res_35_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_18_hi_lo_lo_lo = {wire_res_35_58,wire_res_35_57,wire_res_35_56,wire_res_35_55,wire_res_35_54,
    wire_res_35_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_18_hi_lo_lo = {wire_res_35_65,wire_res_35_64,wire_res_35_63,wire_res_35_62,wire_res_35_61,
    wire_res_35_60,wire_res_35_59,result_reg_w_18_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_18_hi_lo = {wire_res_35_78,wire_res_35_77,wire_res_35_76,wire_res_35_75,wire_res_35_74,
    wire_res_35_73,wire_res_35_72,result_reg_w_18_hi_lo_hi_lo,result_reg_w_18_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_18_hi = {wire_res_35_105,wire_res_35_104,wire_res_35_103,wire_res_35_102,wire_res_35_101,
    wire_res_35_100,wire_res_35_99,result_reg_w_18_hi_hi_hi_lo,result_reg_w_18_hi_hi_lo,result_reg_w_18_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_18_lo_hi_hi_lo = {wire_res_35_45,wire_res_35_44,wire_res_35_43,wire_res_35_42,wire_res_35_41,
    wire_res_35_40,wire_res_35_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_18_lo_hi_lo_lo = {wire_res_35_31,wire_res_35_30,wire_res_35_29,wire_res_35_28,wire_res_35_27,
    wire_res_35_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_18_lo_hi_lo = {wire_res_35_38,wire_res_35_37,wire_res_35_36,wire_res_35_35,wire_res_35_34,
    wire_res_35_33,wire_res_35_32,result_reg_w_18_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_18_lo_lo_hi_lo = {wire_res_35_18,wire_res_35_17,wire_res_35_16,wire_res_35_15,wire_res_35_14,
    wire_res_35_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_18_lo_lo_lo_lo = {wire_res_35_5,wire_res_35_4,wire_res_35_3,wire_res_35_2,wire_res_35_1,
    wire_res_35_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_18_lo_lo_lo = {wire_res_35_12,wire_res_35_11,wire_res_35_10,wire_res_35_9,wire_res_35_8,
    wire_res_35_7,wire_res_35_6,result_reg_w_18_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_18_lo_lo = {wire_res_35_25,wire_res_35_24,wire_res_35_23,wire_res_35_22,wire_res_35_21,
    wire_res_35_20,wire_res_35_19,result_reg_w_18_lo_lo_hi_lo,result_reg_w_18_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_18_lo = {wire_res_35_52,wire_res_35_51,wire_res_35_50,wire_res_35_49,wire_res_35_48,
    wire_res_35_47,wire_res_35_46,result_reg_w_18_lo_hi_hi_lo,result_reg_w_18_lo_hi_lo,result_reg_w_18_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_18 = {result_reg_w_18_hi,result_reg_w_18_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_36_0 = result_reg_w_18[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_1 = result_reg_w_18[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_2 = result_reg_w_18[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_3 = result_reg_w_18[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_4 = result_reg_w_18[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_5 = result_reg_w_18[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_6 = result_reg_w_18[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_7 = result_reg_w_18[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_8 = result_reg_w_18[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_9 = result_reg_w_18[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_10 = result_reg_w_18[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_11 = result_reg_w_18[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_12 = result_reg_w_18[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_13 = result_reg_w_18[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_14 = result_reg_w_18[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_15 = result_reg_w_18[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_16 = result_reg_w_18[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_17 = result_reg_w_18[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_18 = result_reg_w_18[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_19 = result_reg_w_18[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_20 = result_reg_w_18[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_21 = result_reg_w_18[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_22 = result_reg_w_18[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_23 = result_reg_w_18[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_24 = result_reg_w_18[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_25 = result_reg_w_18[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_26 = result_reg_w_18[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_27 = result_reg_w_18[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_28 = result_reg_w_18[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_29 = result_reg_w_18[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_30 = result_reg_w_18[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_31 = result_reg_w_18[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_32 = result_reg_w_18[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_33 = result_reg_w_18[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_34 = result_reg_w_18[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_35 = result_reg_w_18[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_36 = result_reg_w_18[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_37 = result_reg_w_18[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_38 = result_reg_w_18[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_39 = result_reg_w_18[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_40 = result_reg_w_18[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_41 = result_reg_w_18[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_42 = result_reg_w_18[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_43 = result_reg_w_18[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_44 = result_reg_w_18[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_45 = result_reg_w_18[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_46 = result_reg_w_18[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_47 = result_reg_w_18[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_48 = result_reg_w_18[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_49 = result_reg_w_18[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_50 = result_reg_w_18[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_51 = result_reg_w_18[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_52 = result_reg_w_18[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_53 = result_reg_w_18[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_54 = result_reg_w_18[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_55 = result_reg_w_18[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_56 = result_reg_w_18[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_57 = result_reg_w_18[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_58 = result_reg_w_18[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_59 = result_reg_w_18[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_60 = result_reg_w_18[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_61 = result_reg_w_18[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_62 = result_reg_w_18[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_63 = result_reg_w_18[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_64 = result_reg_w_18[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_65 = result_reg_w_18[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_66 = result_reg_w_18[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_67 = result_reg_w_18[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_69 = result_reg_w_18[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_70 = result_reg_w_18[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_71 = result_reg_w_18[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_72 = result_reg_w_18[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_73 = result_reg_w_18[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_74 = result_reg_w_18[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_75 = result_reg_w_18[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_76 = result_reg_w_18[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_77 = result_reg_w_18[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_78 = result_reg_w_18[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_79 = result_reg_w_18[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_80 = result_reg_w_18[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_81 = result_reg_w_18[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_82 = result_reg_w_18[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_83 = result_reg_w_18[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_84 = result_reg_w_18[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_85 = result_reg_w_18[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_86 = result_reg_w_18[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_87 = result_reg_w_18[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_88 = result_reg_w_18[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_89 = result_reg_w_18[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_90 = result_reg_w_18[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_91 = result_reg_w_18[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_92 = result_reg_w_18[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_93 = result_reg_w_18[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_94 = result_reg_w_18[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_95 = result_reg_w_18[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_96 = result_reg_w_18[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_97 = result_reg_w_18[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_98 = result_reg_w_18[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_99 = result_reg_w_18[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_100 = result_reg_w_18[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_101 = result_reg_w_18[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_102 = result_reg_w_18[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_103 = result_reg_w_18[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_104 = result_reg_w_18[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_36_105 = result_reg_w_18[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_0 = result_reg_r_18[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_1 = result_reg_r_18[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_2 = result_reg_r_18[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_3 = result_reg_r_18[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_4 = result_reg_r_18[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_5 = result_reg_r_18[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_6 = result_reg_r_18[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_7 = result_reg_r_18[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_8 = result_reg_r_18[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_9 = result_reg_r_18[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_10 = result_reg_r_18[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_11 = result_reg_r_18[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_12 = result_reg_r_18[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_13 = result_reg_r_18[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_14 = result_reg_r_18[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_15 = result_reg_r_18[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_16 = result_reg_r_18[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_17 = result_reg_r_18[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_18 = result_reg_r_18[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_19 = result_reg_r_18[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_20 = result_reg_r_18[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_21 = result_reg_r_18[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_22 = result_reg_r_18[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_23 = result_reg_r_18[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_24 = result_reg_r_18[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_25 = result_reg_r_18[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_26 = result_reg_r_18[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_27 = result_reg_r_18[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_28 = result_reg_r_18[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_29 = result_reg_r_18[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_30 = result_reg_r_18[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_31 = result_reg_r_18[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_32 = result_reg_r_18[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_33 = result_reg_r_18[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_34 = result_reg_r_18[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_35 = result_reg_r_18[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_36 = result_reg_r_18[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_37 = result_reg_r_18[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_38 = result_reg_r_18[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_39 = result_reg_r_18[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_40 = result_reg_r_18[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_41 = result_reg_r_18[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_42 = result_reg_r_18[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_43 = result_reg_r_18[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_44 = result_reg_r_18[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_45 = result_reg_r_18[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_46 = result_reg_r_18[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_47 = result_reg_r_18[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_48 = result_reg_r_18[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_49 = result_reg_r_18[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_50 = result_reg_r_18[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_51 = result_reg_r_18[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_52 = result_reg_r_18[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_53 = result_reg_r_18[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_54 = result_reg_r_18[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_55 = result_reg_r_18[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_56 = result_reg_r_18[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_57 = result_reg_r_18[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_58 = result_reg_r_18[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_59 = result_reg_r_18[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_60 = result_reg_r_18[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_61 = result_reg_r_18[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_62 = result_reg_r_18[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_63 = result_reg_r_18[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_64 = result_reg_r_18[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_65 = result_reg_r_18[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_66 = result_reg_r_18[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_68 = result_reg_r_18[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_69 = result_reg_r_18[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_70 = result_reg_r_18[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_71 = result_reg_r_18[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_72 = result_reg_r_18[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_73 = result_reg_r_18[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_74 = result_reg_r_18[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_75 = result_reg_r_18[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_76 = result_reg_r_18[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_77 = result_reg_r_18[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_78 = result_reg_r_18[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_79 = result_reg_r_18[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_80 = result_reg_r_18[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_81 = result_reg_r_18[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_82 = result_reg_r_18[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_83 = result_reg_r_18[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_84 = result_reg_r_18[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_85 = result_reg_r_18[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_86 = result_reg_r_18[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_87 = result_reg_r_18[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_88 = result_reg_r_18[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_89 = result_reg_r_18[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_90 = result_reg_r_18[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_91 = result_reg_r_18[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_92 = result_reg_r_18[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_93 = result_reg_r_18[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_94 = result_reg_r_18[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_95 = result_reg_r_18[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_96 = result_reg_r_18[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_97 = result_reg_r_18[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_98 = result_reg_r_18[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_99 = result_reg_r_18[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_100 = result_reg_r_18[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_101 = result_reg_r_18[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_102 = result_reg_r_18[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_103 = result_reg_r_18[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_104 = result_reg_r_18[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_37_105 = result_reg_r_18[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_19_hi_hi_hi_lo = {wire_res_37_98,wire_res_37_97,wire_res_37_96,wire_res_37_95,wire_res_37_94,
    wire_res_37_93,wire_res_37_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_19_hi_hi_lo_lo = {wire_res_37_84,wire_res_37_83,wire_res_37_82,wire_res_37_81,wire_res_37_80,
    wire_res_37_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_19_hi_hi_lo = {wire_res_37_91,wire_res_37_90,wire_res_37_89,wire_res_37_88,wire_res_37_87,
    wire_res_37_86,wire_res_37_85,result_reg_w_19_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [172:0] _T_11312 = {b_aux_reg_r_18, 67'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [172:0] _GEN_1290 = {{67'd0}, a_aux_reg_r_18}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_37_67 = _GEN_1290 >= _T_11312; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_19_hi_lo_hi_lo = {wire_res_37_71,wire_res_37_70,wire_res_37_69,wire_res_37_68,wire_res_37_67,
    wire_res_37_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_19_hi_lo_lo_lo = {wire_res_37_58,wire_res_37_57,wire_res_37_56,wire_res_37_55,wire_res_37_54,
    wire_res_37_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_19_hi_lo_lo = {wire_res_37_65,wire_res_37_64,wire_res_37_63,wire_res_37_62,wire_res_37_61,
    wire_res_37_60,wire_res_37_59,result_reg_w_19_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_19_hi_lo = {wire_res_37_78,wire_res_37_77,wire_res_37_76,wire_res_37_75,wire_res_37_74,
    wire_res_37_73,wire_res_37_72,result_reg_w_19_hi_lo_hi_lo,result_reg_w_19_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_19_hi = {wire_res_37_105,wire_res_37_104,wire_res_37_103,wire_res_37_102,wire_res_37_101,
    wire_res_37_100,wire_res_37_99,result_reg_w_19_hi_hi_hi_lo,result_reg_w_19_hi_hi_lo,result_reg_w_19_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_19_lo_hi_hi_lo = {wire_res_37_45,wire_res_37_44,wire_res_37_43,wire_res_37_42,wire_res_37_41,
    wire_res_37_40,wire_res_37_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_19_lo_hi_lo_lo = {wire_res_37_31,wire_res_37_30,wire_res_37_29,wire_res_37_28,wire_res_37_27,
    wire_res_37_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_19_lo_hi_lo = {wire_res_37_38,wire_res_37_37,wire_res_37_36,wire_res_37_35,wire_res_37_34,
    wire_res_37_33,wire_res_37_32,result_reg_w_19_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_19_lo_lo_hi_lo = {wire_res_37_18,wire_res_37_17,wire_res_37_16,wire_res_37_15,wire_res_37_14,
    wire_res_37_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_19_lo_lo_lo_lo = {wire_res_37_5,wire_res_37_4,wire_res_37_3,wire_res_37_2,wire_res_37_1,
    wire_res_37_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_19_lo_lo_lo = {wire_res_37_12,wire_res_37_11,wire_res_37_10,wire_res_37_9,wire_res_37_8,
    wire_res_37_7,wire_res_37_6,result_reg_w_19_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_19_lo_lo = {wire_res_37_25,wire_res_37_24,wire_res_37_23,wire_res_37_22,wire_res_37_21,
    wire_res_37_20,wire_res_37_19,result_reg_w_19_lo_lo_hi_lo,result_reg_w_19_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_19_lo = {wire_res_37_52,wire_res_37_51,wire_res_37_50,wire_res_37_49,wire_res_37_48,
    wire_res_37_47,wire_res_37_46,result_reg_w_19_lo_hi_hi_lo,result_reg_w_19_lo_hi_lo,result_reg_w_19_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_19 = {result_reg_w_19_hi,result_reg_w_19_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_38_0 = result_reg_w_19[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_1 = result_reg_w_19[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_2 = result_reg_w_19[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_3 = result_reg_w_19[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_4 = result_reg_w_19[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_5 = result_reg_w_19[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_6 = result_reg_w_19[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_7 = result_reg_w_19[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_8 = result_reg_w_19[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_9 = result_reg_w_19[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_10 = result_reg_w_19[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_11 = result_reg_w_19[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_12 = result_reg_w_19[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_13 = result_reg_w_19[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_14 = result_reg_w_19[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_15 = result_reg_w_19[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_16 = result_reg_w_19[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_17 = result_reg_w_19[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_18 = result_reg_w_19[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_19 = result_reg_w_19[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_20 = result_reg_w_19[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_21 = result_reg_w_19[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_22 = result_reg_w_19[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_23 = result_reg_w_19[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_24 = result_reg_w_19[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_25 = result_reg_w_19[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_26 = result_reg_w_19[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_27 = result_reg_w_19[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_28 = result_reg_w_19[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_29 = result_reg_w_19[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_30 = result_reg_w_19[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_31 = result_reg_w_19[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_32 = result_reg_w_19[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_33 = result_reg_w_19[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_34 = result_reg_w_19[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_35 = result_reg_w_19[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_36 = result_reg_w_19[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_37 = result_reg_w_19[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_38 = result_reg_w_19[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_39 = result_reg_w_19[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_40 = result_reg_w_19[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_41 = result_reg_w_19[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_42 = result_reg_w_19[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_43 = result_reg_w_19[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_44 = result_reg_w_19[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_45 = result_reg_w_19[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_46 = result_reg_w_19[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_47 = result_reg_w_19[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_48 = result_reg_w_19[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_49 = result_reg_w_19[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_50 = result_reg_w_19[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_51 = result_reg_w_19[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_52 = result_reg_w_19[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_53 = result_reg_w_19[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_54 = result_reg_w_19[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_55 = result_reg_w_19[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_56 = result_reg_w_19[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_57 = result_reg_w_19[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_58 = result_reg_w_19[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_59 = result_reg_w_19[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_60 = result_reg_w_19[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_61 = result_reg_w_19[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_62 = result_reg_w_19[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_63 = result_reg_w_19[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_64 = result_reg_w_19[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_65 = result_reg_w_19[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_67 = result_reg_w_19[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_68 = result_reg_w_19[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_69 = result_reg_w_19[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_70 = result_reg_w_19[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_71 = result_reg_w_19[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_72 = result_reg_w_19[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_73 = result_reg_w_19[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_74 = result_reg_w_19[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_75 = result_reg_w_19[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_76 = result_reg_w_19[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_77 = result_reg_w_19[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_78 = result_reg_w_19[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_79 = result_reg_w_19[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_80 = result_reg_w_19[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_81 = result_reg_w_19[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_82 = result_reg_w_19[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_83 = result_reg_w_19[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_84 = result_reg_w_19[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_85 = result_reg_w_19[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_86 = result_reg_w_19[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_87 = result_reg_w_19[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_88 = result_reg_w_19[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_89 = result_reg_w_19[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_90 = result_reg_w_19[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_91 = result_reg_w_19[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_92 = result_reg_w_19[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_93 = result_reg_w_19[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_94 = result_reg_w_19[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_95 = result_reg_w_19[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_96 = result_reg_w_19[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_97 = result_reg_w_19[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_98 = result_reg_w_19[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_99 = result_reg_w_19[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_100 = result_reg_w_19[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_101 = result_reg_w_19[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_102 = result_reg_w_19[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_103 = result_reg_w_19[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_104 = result_reg_w_19[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_38_105 = result_reg_w_19[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_0 = result_reg_r_19[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_1 = result_reg_r_19[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_2 = result_reg_r_19[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_3 = result_reg_r_19[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_4 = result_reg_r_19[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_5 = result_reg_r_19[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_6 = result_reg_r_19[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_7 = result_reg_r_19[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_8 = result_reg_r_19[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_9 = result_reg_r_19[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_10 = result_reg_r_19[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_11 = result_reg_r_19[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_12 = result_reg_r_19[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_13 = result_reg_r_19[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_14 = result_reg_r_19[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_15 = result_reg_r_19[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_16 = result_reg_r_19[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_17 = result_reg_r_19[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_18 = result_reg_r_19[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_19 = result_reg_r_19[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_20 = result_reg_r_19[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_21 = result_reg_r_19[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_22 = result_reg_r_19[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_23 = result_reg_r_19[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_24 = result_reg_r_19[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_25 = result_reg_r_19[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_26 = result_reg_r_19[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_27 = result_reg_r_19[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_28 = result_reg_r_19[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_29 = result_reg_r_19[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_30 = result_reg_r_19[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_31 = result_reg_r_19[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_32 = result_reg_r_19[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_33 = result_reg_r_19[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_34 = result_reg_r_19[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_35 = result_reg_r_19[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_36 = result_reg_r_19[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_37 = result_reg_r_19[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_38 = result_reg_r_19[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_39 = result_reg_r_19[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_40 = result_reg_r_19[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_41 = result_reg_r_19[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_42 = result_reg_r_19[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_43 = result_reg_r_19[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_44 = result_reg_r_19[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_45 = result_reg_r_19[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_46 = result_reg_r_19[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_47 = result_reg_r_19[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_48 = result_reg_r_19[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_49 = result_reg_r_19[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_50 = result_reg_r_19[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_51 = result_reg_r_19[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_52 = result_reg_r_19[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_53 = result_reg_r_19[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_54 = result_reg_r_19[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_55 = result_reg_r_19[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_56 = result_reg_r_19[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_57 = result_reg_r_19[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_58 = result_reg_r_19[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_59 = result_reg_r_19[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_60 = result_reg_r_19[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_61 = result_reg_r_19[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_62 = result_reg_r_19[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_63 = result_reg_r_19[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_64 = result_reg_r_19[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_66 = result_reg_r_19[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_67 = result_reg_r_19[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_68 = result_reg_r_19[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_69 = result_reg_r_19[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_70 = result_reg_r_19[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_71 = result_reg_r_19[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_72 = result_reg_r_19[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_73 = result_reg_r_19[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_74 = result_reg_r_19[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_75 = result_reg_r_19[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_76 = result_reg_r_19[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_77 = result_reg_r_19[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_78 = result_reg_r_19[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_79 = result_reg_r_19[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_80 = result_reg_r_19[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_81 = result_reg_r_19[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_82 = result_reg_r_19[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_83 = result_reg_r_19[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_84 = result_reg_r_19[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_85 = result_reg_r_19[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_86 = result_reg_r_19[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_87 = result_reg_r_19[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_88 = result_reg_r_19[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_89 = result_reg_r_19[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_90 = result_reg_r_19[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_91 = result_reg_r_19[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_92 = result_reg_r_19[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_93 = result_reg_r_19[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_94 = result_reg_r_19[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_95 = result_reg_r_19[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_96 = result_reg_r_19[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_97 = result_reg_r_19[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_98 = result_reg_r_19[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_99 = result_reg_r_19[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_100 = result_reg_r_19[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_101 = result_reg_r_19[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_102 = result_reg_r_19[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_103 = result_reg_r_19[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_104 = result_reg_r_19[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_39_105 = result_reg_r_19[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_20_hi_hi_hi_lo = {wire_res_39_98,wire_res_39_97,wire_res_39_96,wire_res_39_95,wire_res_39_94,
    wire_res_39_93,wire_res_39_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_20_hi_hi_lo_lo = {wire_res_39_84,wire_res_39_83,wire_res_39_82,wire_res_39_81,wire_res_39_80,
    wire_res_39_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_20_hi_hi_lo = {wire_res_39_91,wire_res_39_90,wire_res_39_89,wire_res_39_88,wire_res_39_87,
    wire_res_39_86,wire_res_39_85,result_reg_w_20_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_20_hi_lo_hi_lo = {wire_res_39_71,wire_res_39_70,wire_res_39_69,wire_res_39_68,wire_res_39_67,
    wire_res_39_66}; // @[BinaryDesigns2.scala 231:46]
  wire [170:0] _T_11316 = {b_aux_reg_r_19, 65'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [170:0] _GEN_1291 = {{65'd0}, a_aux_reg_r_19}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_39_65 = _GEN_1291 >= _T_11316; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_20_hi_lo_lo_lo = {wire_res_39_58,wire_res_39_57,wire_res_39_56,wire_res_39_55,wire_res_39_54,
    wire_res_39_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_20_hi_lo_lo = {wire_res_39_65,wire_res_39_64,wire_res_39_63,wire_res_39_62,wire_res_39_61,
    wire_res_39_60,wire_res_39_59,result_reg_w_20_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_20_hi_lo = {wire_res_39_78,wire_res_39_77,wire_res_39_76,wire_res_39_75,wire_res_39_74,
    wire_res_39_73,wire_res_39_72,result_reg_w_20_hi_lo_hi_lo,result_reg_w_20_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_20_hi = {wire_res_39_105,wire_res_39_104,wire_res_39_103,wire_res_39_102,wire_res_39_101,
    wire_res_39_100,wire_res_39_99,result_reg_w_20_hi_hi_hi_lo,result_reg_w_20_hi_hi_lo,result_reg_w_20_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_20_lo_hi_hi_lo = {wire_res_39_45,wire_res_39_44,wire_res_39_43,wire_res_39_42,wire_res_39_41,
    wire_res_39_40,wire_res_39_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_20_lo_hi_lo_lo = {wire_res_39_31,wire_res_39_30,wire_res_39_29,wire_res_39_28,wire_res_39_27,
    wire_res_39_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_20_lo_hi_lo = {wire_res_39_38,wire_res_39_37,wire_res_39_36,wire_res_39_35,wire_res_39_34,
    wire_res_39_33,wire_res_39_32,result_reg_w_20_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_20_lo_lo_hi_lo = {wire_res_39_18,wire_res_39_17,wire_res_39_16,wire_res_39_15,wire_res_39_14,
    wire_res_39_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_20_lo_lo_lo_lo = {wire_res_39_5,wire_res_39_4,wire_res_39_3,wire_res_39_2,wire_res_39_1,
    wire_res_39_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_20_lo_lo_lo = {wire_res_39_12,wire_res_39_11,wire_res_39_10,wire_res_39_9,wire_res_39_8,
    wire_res_39_7,wire_res_39_6,result_reg_w_20_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_20_lo_lo = {wire_res_39_25,wire_res_39_24,wire_res_39_23,wire_res_39_22,wire_res_39_21,
    wire_res_39_20,wire_res_39_19,result_reg_w_20_lo_lo_hi_lo,result_reg_w_20_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_20_lo = {wire_res_39_52,wire_res_39_51,wire_res_39_50,wire_res_39_49,wire_res_39_48,
    wire_res_39_47,wire_res_39_46,result_reg_w_20_lo_hi_hi_lo,result_reg_w_20_lo_hi_lo,result_reg_w_20_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_20 = {result_reg_w_20_hi,result_reg_w_20_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_40_0 = result_reg_w_20[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_1 = result_reg_w_20[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_2 = result_reg_w_20[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_3 = result_reg_w_20[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_4 = result_reg_w_20[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_5 = result_reg_w_20[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_6 = result_reg_w_20[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_7 = result_reg_w_20[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_8 = result_reg_w_20[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_9 = result_reg_w_20[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_10 = result_reg_w_20[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_11 = result_reg_w_20[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_12 = result_reg_w_20[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_13 = result_reg_w_20[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_14 = result_reg_w_20[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_15 = result_reg_w_20[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_16 = result_reg_w_20[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_17 = result_reg_w_20[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_18 = result_reg_w_20[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_19 = result_reg_w_20[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_20 = result_reg_w_20[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_21 = result_reg_w_20[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_22 = result_reg_w_20[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_23 = result_reg_w_20[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_24 = result_reg_w_20[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_25 = result_reg_w_20[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_26 = result_reg_w_20[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_27 = result_reg_w_20[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_28 = result_reg_w_20[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_29 = result_reg_w_20[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_30 = result_reg_w_20[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_31 = result_reg_w_20[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_32 = result_reg_w_20[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_33 = result_reg_w_20[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_34 = result_reg_w_20[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_35 = result_reg_w_20[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_36 = result_reg_w_20[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_37 = result_reg_w_20[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_38 = result_reg_w_20[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_39 = result_reg_w_20[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_40 = result_reg_w_20[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_41 = result_reg_w_20[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_42 = result_reg_w_20[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_43 = result_reg_w_20[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_44 = result_reg_w_20[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_45 = result_reg_w_20[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_46 = result_reg_w_20[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_47 = result_reg_w_20[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_48 = result_reg_w_20[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_49 = result_reg_w_20[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_50 = result_reg_w_20[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_51 = result_reg_w_20[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_52 = result_reg_w_20[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_53 = result_reg_w_20[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_54 = result_reg_w_20[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_55 = result_reg_w_20[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_56 = result_reg_w_20[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_57 = result_reg_w_20[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_58 = result_reg_w_20[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_59 = result_reg_w_20[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_60 = result_reg_w_20[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_61 = result_reg_w_20[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_62 = result_reg_w_20[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_63 = result_reg_w_20[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_65 = result_reg_w_20[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_66 = result_reg_w_20[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_67 = result_reg_w_20[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_68 = result_reg_w_20[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_69 = result_reg_w_20[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_70 = result_reg_w_20[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_71 = result_reg_w_20[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_72 = result_reg_w_20[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_73 = result_reg_w_20[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_74 = result_reg_w_20[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_75 = result_reg_w_20[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_76 = result_reg_w_20[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_77 = result_reg_w_20[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_78 = result_reg_w_20[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_79 = result_reg_w_20[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_80 = result_reg_w_20[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_81 = result_reg_w_20[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_82 = result_reg_w_20[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_83 = result_reg_w_20[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_84 = result_reg_w_20[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_85 = result_reg_w_20[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_86 = result_reg_w_20[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_87 = result_reg_w_20[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_88 = result_reg_w_20[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_89 = result_reg_w_20[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_90 = result_reg_w_20[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_91 = result_reg_w_20[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_92 = result_reg_w_20[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_93 = result_reg_w_20[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_94 = result_reg_w_20[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_95 = result_reg_w_20[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_96 = result_reg_w_20[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_97 = result_reg_w_20[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_98 = result_reg_w_20[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_99 = result_reg_w_20[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_100 = result_reg_w_20[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_101 = result_reg_w_20[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_102 = result_reg_w_20[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_103 = result_reg_w_20[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_104 = result_reg_w_20[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_40_105 = result_reg_w_20[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_0 = result_reg_r_20[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_1 = result_reg_r_20[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_2 = result_reg_r_20[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_3 = result_reg_r_20[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_4 = result_reg_r_20[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_5 = result_reg_r_20[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_6 = result_reg_r_20[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_7 = result_reg_r_20[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_8 = result_reg_r_20[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_9 = result_reg_r_20[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_10 = result_reg_r_20[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_11 = result_reg_r_20[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_12 = result_reg_r_20[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_13 = result_reg_r_20[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_14 = result_reg_r_20[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_15 = result_reg_r_20[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_16 = result_reg_r_20[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_17 = result_reg_r_20[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_18 = result_reg_r_20[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_19 = result_reg_r_20[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_20 = result_reg_r_20[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_21 = result_reg_r_20[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_22 = result_reg_r_20[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_23 = result_reg_r_20[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_24 = result_reg_r_20[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_25 = result_reg_r_20[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_26 = result_reg_r_20[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_27 = result_reg_r_20[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_28 = result_reg_r_20[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_29 = result_reg_r_20[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_30 = result_reg_r_20[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_31 = result_reg_r_20[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_32 = result_reg_r_20[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_33 = result_reg_r_20[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_34 = result_reg_r_20[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_35 = result_reg_r_20[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_36 = result_reg_r_20[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_37 = result_reg_r_20[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_38 = result_reg_r_20[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_39 = result_reg_r_20[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_40 = result_reg_r_20[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_41 = result_reg_r_20[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_42 = result_reg_r_20[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_43 = result_reg_r_20[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_44 = result_reg_r_20[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_45 = result_reg_r_20[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_46 = result_reg_r_20[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_47 = result_reg_r_20[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_48 = result_reg_r_20[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_49 = result_reg_r_20[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_50 = result_reg_r_20[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_51 = result_reg_r_20[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_52 = result_reg_r_20[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_53 = result_reg_r_20[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_54 = result_reg_r_20[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_55 = result_reg_r_20[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_56 = result_reg_r_20[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_57 = result_reg_r_20[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_58 = result_reg_r_20[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_59 = result_reg_r_20[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_60 = result_reg_r_20[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_61 = result_reg_r_20[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_62 = result_reg_r_20[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_64 = result_reg_r_20[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_65 = result_reg_r_20[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_66 = result_reg_r_20[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_67 = result_reg_r_20[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_68 = result_reg_r_20[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_69 = result_reg_r_20[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_70 = result_reg_r_20[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_71 = result_reg_r_20[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_72 = result_reg_r_20[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_73 = result_reg_r_20[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_74 = result_reg_r_20[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_75 = result_reg_r_20[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_76 = result_reg_r_20[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_77 = result_reg_r_20[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_78 = result_reg_r_20[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_79 = result_reg_r_20[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_80 = result_reg_r_20[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_81 = result_reg_r_20[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_82 = result_reg_r_20[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_83 = result_reg_r_20[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_84 = result_reg_r_20[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_85 = result_reg_r_20[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_86 = result_reg_r_20[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_87 = result_reg_r_20[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_88 = result_reg_r_20[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_89 = result_reg_r_20[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_90 = result_reg_r_20[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_91 = result_reg_r_20[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_92 = result_reg_r_20[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_93 = result_reg_r_20[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_94 = result_reg_r_20[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_95 = result_reg_r_20[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_96 = result_reg_r_20[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_97 = result_reg_r_20[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_98 = result_reg_r_20[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_99 = result_reg_r_20[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_100 = result_reg_r_20[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_101 = result_reg_r_20[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_102 = result_reg_r_20[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_103 = result_reg_r_20[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_104 = result_reg_r_20[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_41_105 = result_reg_r_20[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_21_hi_hi_hi_lo = {wire_res_41_98,wire_res_41_97,wire_res_41_96,wire_res_41_95,wire_res_41_94,
    wire_res_41_93,wire_res_41_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_21_hi_hi_lo_lo = {wire_res_41_84,wire_res_41_83,wire_res_41_82,wire_res_41_81,wire_res_41_80,
    wire_res_41_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_21_hi_hi_lo = {wire_res_41_91,wire_res_41_90,wire_res_41_89,wire_res_41_88,wire_res_41_87,
    wire_res_41_86,wire_res_41_85,result_reg_w_21_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_21_hi_lo_hi_lo = {wire_res_41_71,wire_res_41_70,wire_res_41_69,wire_res_41_68,wire_res_41_67,
    wire_res_41_66}; // @[BinaryDesigns2.scala 231:46]
  wire [168:0] _T_11320 = {b_aux_reg_r_20, 63'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [168:0] _GEN_1292 = {{63'd0}, a_aux_reg_r_20}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_41_63 = _GEN_1292 >= _T_11320; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_21_hi_lo_lo_lo = {wire_res_41_58,wire_res_41_57,wire_res_41_56,wire_res_41_55,wire_res_41_54,
    wire_res_41_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_21_hi_lo_lo = {wire_res_41_65,wire_res_41_64,wire_res_41_63,wire_res_41_62,wire_res_41_61,
    wire_res_41_60,wire_res_41_59,result_reg_w_21_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_21_hi_lo = {wire_res_41_78,wire_res_41_77,wire_res_41_76,wire_res_41_75,wire_res_41_74,
    wire_res_41_73,wire_res_41_72,result_reg_w_21_hi_lo_hi_lo,result_reg_w_21_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_21_hi = {wire_res_41_105,wire_res_41_104,wire_res_41_103,wire_res_41_102,wire_res_41_101,
    wire_res_41_100,wire_res_41_99,result_reg_w_21_hi_hi_hi_lo,result_reg_w_21_hi_hi_lo,result_reg_w_21_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_21_lo_hi_hi_lo = {wire_res_41_45,wire_res_41_44,wire_res_41_43,wire_res_41_42,wire_res_41_41,
    wire_res_41_40,wire_res_41_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_21_lo_hi_lo_lo = {wire_res_41_31,wire_res_41_30,wire_res_41_29,wire_res_41_28,wire_res_41_27,
    wire_res_41_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_21_lo_hi_lo = {wire_res_41_38,wire_res_41_37,wire_res_41_36,wire_res_41_35,wire_res_41_34,
    wire_res_41_33,wire_res_41_32,result_reg_w_21_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_21_lo_lo_hi_lo = {wire_res_41_18,wire_res_41_17,wire_res_41_16,wire_res_41_15,wire_res_41_14,
    wire_res_41_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_21_lo_lo_lo_lo = {wire_res_41_5,wire_res_41_4,wire_res_41_3,wire_res_41_2,wire_res_41_1,
    wire_res_41_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_21_lo_lo_lo = {wire_res_41_12,wire_res_41_11,wire_res_41_10,wire_res_41_9,wire_res_41_8,
    wire_res_41_7,wire_res_41_6,result_reg_w_21_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_21_lo_lo = {wire_res_41_25,wire_res_41_24,wire_res_41_23,wire_res_41_22,wire_res_41_21,
    wire_res_41_20,wire_res_41_19,result_reg_w_21_lo_lo_hi_lo,result_reg_w_21_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_21_lo = {wire_res_41_52,wire_res_41_51,wire_res_41_50,wire_res_41_49,wire_res_41_48,
    wire_res_41_47,wire_res_41_46,result_reg_w_21_lo_hi_hi_lo,result_reg_w_21_lo_hi_lo,result_reg_w_21_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_21 = {result_reg_w_21_hi,result_reg_w_21_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_42_0 = result_reg_w_21[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_1 = result_reg_w_21[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_2 = result_reg_w_21[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_3 = result_reg_w_21[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_4 = result_reg_w_21[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_5 = result_reg_w_21[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_6 = result_reg_w_21[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_7 = result_reg_w_21[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_8 = result_reg_w_21[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_9 = result_reg_w_21[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_10 = result_reg_w_21[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_11 = result_reg_w_21[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_12 = result_reg_w_21[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_13 = result_reg_w_21[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_14 = result_reg_w_21[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_15 = result_reg_w_21[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_16 = result_reg_w_21[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_17 = result_reg_w_21[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_18 = result_reg_w_21[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_19 = result_reg_w_21[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_20 = result_reg_w_21[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_21 = result_reg_w_21[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_22 = result_reg_w_21[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_23 = result_reg_w_21[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_24 = result_reg_w_21[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_25 = result_reg_w_21[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_26 = result_reg_w_21[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_27 = result_reg_w_21[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_28 = result_reg_w_21[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_29 = result_reg_w_21[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_30 = result_reg_w_21[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_31 = result_reg_w_21[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_32 = result_reg_w_21[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_33 = result_reg_w_21[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_34 = result_reg_w_21[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_35 = result_reg_w_21[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_36 = result_reg_w_21[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_37 = result_reg_w_21[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_38 = result_reg_w_21[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_39 = result_reg_w_21[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_40 = result_reg_w_21[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_41 = result_reg_w_21[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_42 = result_reg_w_21[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_43 = result_reg_w_21[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_44 = result_reg_w_21[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_45 = result_reg_w_21[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_46 = result_reg_w_21[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_47 = result_reg_w_21[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_48 = result_reg_w_21[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_49 = result_reg_w_21[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_50 = result_reg_w_21[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_51 = result_reg_w_21[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_52 = result_reg_w_21[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_53 = result_reg_w_21[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_54 = result_reg_w_21[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_55 = result_reg_w_21[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_56 = result_reg_w_21[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_57 = result_reg_w_21[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_58 = result_reg_w_21[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_59 = result_reg_w_21[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_60 = result_reg_w_21[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_61 = result_reg_w_21[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_63 = result_reg_w_21[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_64 = result_reg_w_21[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_65 = result_reg_w_21[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_66 = result_reg_w_21[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_67 = result_reg_w_21[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_68 = result_reg_w_21[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_69 = result_reg_w_21[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_70 = result_reg_w_21[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_71 = result_reg_w_21[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_72 = result_reg_w_21[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_73 = result_reg_w_21[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_74 = result_reg_w_21[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_75 = result_reg_w_21[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_76 = result_reg_w_21[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_77 = result_reg_w_21[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_78 = result_reg_w_21[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_79 = result_reg_w_21[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_80 = result_reg_w_21[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_81 = result_reg_w_21[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_82 = result_reg_w_21[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_83 = result_reg_w_21[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_84 = result_reg_w_21[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_85 = result_reg_w_21[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_86 = result_reg_w_21[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_87 = result_reg_w_21[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_88 = result_reg_w_21[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_89 = result_reg_w_21[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_90 = result_reg_w_21[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_91 = result_reg_w_21[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_92 = result_reg_w_21[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_93 = result_reg_w_21[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_94 = result_reg_w_21[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_95 = result_reg_w_21[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_96 = result_reg_w_21[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_97 = result_reg_w_21[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_98 = result_reg_w_21[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_99 = result_reg_w_21[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_100 = result_reg_w_21[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_101 = result_reg_w_21[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_102 = result_reg_w_21[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_103 = result_reg_w_21[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_104 = result_reg_w_21[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_42_105 = result_reg_w_21[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_0 = result_reg_r_21[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_1 = result_reg_r_21[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_2 = result_reg_r_21[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_3 = result_reg_r_21[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_4 = result_reg_r_21[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_5 = result_reg_r_21[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_6 = result_reg_r_21[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_7 = result_reg_r_21[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_8 = result_reg_r_21[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_9 = result_reg_r_21[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_10 = result_reg_r_21[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_11 = result_reg_r_21[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_12 = result_reg_r_21[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_13 = result_reg_r_21[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_14 = result_reg_r_21[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_15 = result_reg_r_21[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_16 = result_reg_r_21[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_17 = result_reg_r_21[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_18 = result_reg_r_21[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_19 = result_reg_r_21[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_20 = result_reg_r_21[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_21 = result_reg_r_21[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_22 = result_reg_r_21[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_23 = result_reg_r_21[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_24 = result_reg_r_21[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_25 = result_reg_r_21[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_26 = result_reg_r_21[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_27 = result_reg_r_21[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_28 = result_reg_r_21[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_29 = result_reg_r_21[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_30 = result_reg_r_21[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_31 = result_reg_r_21[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_32 = result_reg_r_21[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_33 = result_reg_r_21[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_34 = result_reg_r_21[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_35 = result_reg_r_21[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_36 = result_reg_r_21[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_37 = result_reg_r_21[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_38 = result_reg_r_21[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_39 = result_reg_r_21[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_40 = result_reg_r_21[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_41 = result_reg_r_21[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_42 = result_reg_r_21[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_43 = result_reg_r_21[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_44 = result_reg_r_21[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_45 = result_reg_r_21[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_46 = result_reg_r_21[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_47 = result_reg_r_21[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_48 = result_reg_r_21[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_49 = result_reg_r_21[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_50 = result_reg_r_21[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_51 = result_reg_r_21[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_52 = result_reg_r_21[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_53 = result_reg_r_21[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_54 = result_reg_r_21[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_55 = result_reg_r_21[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_56 = result_reg_r_21[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_57 = result_reg_r_21[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_58 = result_reg_r_21[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_59 = result_reg_r_21[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_60 = result_reg_r_21[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_62 = result_reg_r_21[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_63 = result_reg_r_21[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_64 = result_reg_r_21[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_65 = result_reg_r_21[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_66 = result_reg_r_21[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_67 = result_reg_r_21[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_68 = result_reg_r_21[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_69 = result_reg_r_21[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_70 = result_reg_r_21[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_71 = result_reg_r_21[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_72 = result_reg_r_21[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_73 = result_reg_r_21[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_74 = result_reg_r_21[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_75 = result_reg_r_21[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_76 = result_reg_r_21[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_77 = result_reg_r_21[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_78 = result_reg_r_21[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_79 = result_reg_r_21[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_80 = result_reg_r_21[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_81 = result_reg_r_21[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_82 = result_reg_r_21[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_83 = result_reg_r_21[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_84 = result_reg_r_21[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_85 = result_reg_r_21[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_86 = result_reg_r_21[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_87 = result_reg_r_21[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_88 = result_reg_r_21[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_89 = result_reg_r_21[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_90 = result_reg_r_21[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_91 = result_reg_r_21[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_92 = result_reg_r_21[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_93 = result_reg_r_21[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_94 = result_reg_r_21[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_95 = result_reg_r_21[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_96 = result_reg_r_21[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_97 = result_reg_r_21[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_98 = result_reg_r_21[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_99 = result_reg_r_21[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_100 = result_reg_r_21[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_101 = result_reg_r_21[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_102 = result_reg_r_21[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_103 = result_reg_r_21[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_104 = result_reg_r_21[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_43_105 = result_reg_r_21[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_22_hi_hi_hi_lo = {wire_res_43_98,wire_res_43_97,wire_res_43_96,wire_res_43_95,wire_res_43_94,
    wire_res_43_93,wire_res_43_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_22_hi_hi_lo_lo = {wire_res_43_84,wire_res_43_83,wire_res_43_82,wire_res_43_81,wire_res_43_80,
    wire_res_43_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_22_hi_hi_lo = {wire_res_43_91,wire_res_43_90,wire_res_43_89,wire_res_43_88,wire_res_43_87,
    wire_res_43_86,wire_res_43_85,result_reg_w_22_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_22_hi_lo_hi_lo = {wire_res_43_71,wire_res_43_70,wire_res_43_69,wire_res_43_68,wire_res_43_67,
    wire_res_43_66}; // @[BinaryDesigns2.scala 231:46]
  wire [166:0] _T_11324 = {b_aux_reg_r_21, 61'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [166:0] _GEN_1293 = {{61'd0}, a_aux_reg_r_21}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_43_61 = _GEN_1293 >= _T_11324; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_22_hi_lo_lo_lo = {wire_res_43_58,wire_res_43_57,wire_res_43_56,wire_res_43_55,wire_res_43_54,
    wire_res_43_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_22_hi_lo_lo = {wire_res_43_65,wire_res_43_64,wire_res_43_63,wire_res_43_62,wire_res_43_61,
    wire_res_43_60,wire_res_43_59,result_reg_w_22_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_22_hi_lo = {wire_res_43_78,wire_res_43_77,wire_res_43_76,wire_res_43_75,wire_res_43_74,
    wire_res_43_73,wire_res_43_72,result_reg_w_22_hi_lo_hi_lo,result_reg_w_22_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_22_hi = {wire_res_43_105,wire_res_43_104,wire_res_43_103,wire_res_43_102,wire_res_43_101,
    wire_res_43_100,wire_res_43_99,result_reg_w_22_hi_hi_hi_lo,result_reg_w_22_hi_hi_lo,result_reg_w_22_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_22_lo_hi_hi_lo = {wire_res_43_45,wire_res_43_44,wire_res_43_43,wire_res_43_42,wire_res_43_41,
    wire_res_43_40,wire_res_43_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_22_lo_hi_lo_lo = {wire_res_43_31,wire_res_43_30,wire_res_43_29,wire_res_43_28,wire_res_43_27,
    wire_res_43_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_22_lo_hi_lo = {wire_res_43_38,wire_res_43_37,wire_res_43_36,wire_res_43_35,wire_res_43_34,
    wire_res_43_33,wire_res_43_32,result_reg_w_22_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_22_lo_lo_hi_lo = {wire_res_43_18,wire_res_43_17,wire_res_43_16,wire_res_43_15,wire_res_43_14,
    wire_res_43_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_22_lo_lo_lo_lo = {wire_res_43_5,wire_res_43_4,wire_res_43_3,wire_res_43_2,wire_res_43_1,
    wire_res_43_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_22_lo_lo_lo = {wire_res_43_12,wire_res_43_11,wire_res_43_10,wire_res_43_9,wire_res_43_8,
    wire_res_43_7,wire_res_43_6,result_reg_w_22_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_22_lo_lo = {wire_res_43_25,wire_res_43_24,wire_res_43_23,wire_res_43_22,wire_res_43_21,
    wire_res_43_20,wire_res_43_19,result_reg_w_22_lo_lo_hi_lo,result_reg_w_22_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_22_lo = {wire_res_43_52,wire_res_43_51,wire_res_43_50,wire_res_43_49,wire_res_43_48,
    wire_res_43_47,wire_res_43_46,result_reg_w_22_lo_hi_hi_lo,result_reg_w_22_lo_hi_lo,result_reg_w_22_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_22 = {result_reg_w_22_hi,result_reg_w_22_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_44_0 = result_reg_w_22[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_1 = result_reg_w_22[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_2 = result_reg_w_22[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_3 = result_reg_w_22[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_4 = result_reg_w_22[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_5 = result_reg_w_22[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_6 = result_reg_w_22[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_7 = result_reg_w_22[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_8 = result_reg_w_22[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_9 = result_reg_w_22[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_10 = result_reg_w_22[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_11 = result_reg_w_22[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_12 = result_reg_w_22[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_13 = result_reg_w_22[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_14 = result_reg_w_22[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_15 = result_reg_w_22[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_16 = result_reg_w_22[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_17 = result_reg_w_22[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_18 = result_reg_w_22[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_19 = result_reg_w_22[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_20 = result_reg_w_22[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_21 = result_reg_w_22[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_22 = result_reg_w_22[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_23 = result_reg_w_22[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_24 = result_reg_w_22[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_25 = result_reg_w_22[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_26 = result_reg_w_22[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_27 = result_reg_w_22[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_28 = result_reg_w_22[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_29 = result_reg_w_22[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_30 = result_reg_w_22[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_31 = result_reg_w_22[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_32 = result_reg_w_22[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_33 = result_reg_w_22[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_34 = result_reg_w_22[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_35 = result_reg_w_22[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_36 = result_reg_w_22[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_37 = result_reg_w_22[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_38 = result_reg_w_22[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_39 = result_reg_w_22[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_40 = result_reg_w_22[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_41 = result_reg_w_22[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_42 = result_reg_w_22[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_43 = result_reg_w_22[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_44 = result_reg_w_22[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_45 = result_reg_w_22[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_46 = result_reg_w_22[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_47 = result_reg_w_22[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_48 = result_reg_w_22[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_49 = result_reg_w_22[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_50 = result_reg_w_22[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_51 = result_reg_w_22[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_52 = result_reg_w_22[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_53 = result_reg_w_22[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_54 = result_reg_w_22[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_55 = result_reg_w_22[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_56 = result_reg_w_22[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_57 = result_reg_w_22[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_58 = result_reg_w_22[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_59 = result_reg_w_22[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_61 = result_reg_w_22[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_62 = result_reg_w_22[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_63 = result_reg_w_22[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_64 = result_reg_w_22[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_65 = result_reg_w_22[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_66 = result_reg_w_22[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_67 = result_reg_w_22[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_68 = result_reg_w_22[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_69 = result_reg_w_22[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_70 = result_reg_w_22[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_71 = result_reg_w_22[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_72 = result_reg_w_22[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_73 = result_reg_w_22[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_74 = result_reg_w_22[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_75 = result_reg_w_22[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_76 = result_reg_w_22[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_77 = result_reg_w_22[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_78 = result_reg_w_22[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_79 = result_reg_w_22[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_80 = result_reg_w_22[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_81 = result_reg_w_22[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_82 = result_reg_w_22[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_83 = result_reg_w_22[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_84 = result_reg_w_22[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_85 = result_reg_w_22[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_86 = result_reg_w_22[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_87 = result_reg_w_22[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_88 = result_reg_w_22[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_89 = result_reg_w_22[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_90 = result_reg_w_22[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_91 = result_reg_w_22[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_92 = result_reg_w_22[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_93 = result_reg_w_22[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_94 = result_reg_w_22[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_95 = result_reg_w_22[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_96 = result_reg_w_22[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_97 = result_reg_w_22[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_98 = result_reg_w_22[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_99 = result_reg_w_22[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_100 = result_reg_w_22[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_101 = result_reg_w_22[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_102 = result_reg_w_22[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_103 = result_reg_w_22[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_104 = result_reg_w_22[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_44_105 = result_reg_w_22[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_0 = result_reg_r_22[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_1 = result_reg_r_22[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_2 = result_reg_r_22[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_3 = result_reg_r_22[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_4 = result_reg_r_22[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_5 = result_reg_r_22[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_6 = result_reg_r_22[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_7 = result_reg_r_22[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_8 = result_reg_r_22[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_9 = result_reg_r_22[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_10 = result_reg_r_22[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_11 = result_reg_r_22[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_12 = result_reg_r_22[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_13 = result_reg_r_22[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_14 = result_reg_r_22[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_15 = result_reg_r_22[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_16 = result_reg_r_22[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_17 = result_reg_r_22[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_18 = result_reg_r_22[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_19 = result_reg_r_22[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_20 = result_reg_r_22[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_21 = result_reg_r_22[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_22 = result_reg_r_22[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_23 = result_reg_r_22[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_24 = result_reg_r_22[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_25 = result_reg_r_22[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_26 = result_reg_r_22[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_27 = result_reg_r_22[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_28 = result_reg_r_22[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_29 = result_reg_r_22[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_30 = result_reg_r_22[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_31 = result_reg_r_22[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_32 = result_reg_r_22[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_33 = result_reg_r_22[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_34 = result_reg_r_22[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_35 = result_reg_r_22[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_36 = result_reg_r_22[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_37 = result_reg_r_22[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_38 = result_reg_r_22[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_39 = result_reg_r_22[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_40 = result_reg_r_22[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_41 = result_reg_r_22[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_42 = result_reg_r_22[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_43 = result_reg_r_22[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_44 = result_reg_r_22[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_45 = result_reg_r_22[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_46 = result_reg_r_22[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_47 = result_reg_r_22[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_48 = result_reg_r_22[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_49 = result_reg_r_22[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_50 = result_reg_r_22[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_51 = result_reg_r_22[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_52 = result_reg_r_22[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_53 = result_reg_r_22[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_54 = result_reg_r_22[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_55 = result_reg_r_22[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_56 = result_reg_r_22[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_57 = result_reg_r_22[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_58 = result_reg_r_22[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_60 = result_reg_r_22[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_61 = result_reg_r_22[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_62 = result_reg_r_22[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_63 = result_reg_r_22[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_64 = result_reg_r_22[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_65 = result_reg_r_22[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_66 = result_reg_r_22[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_67 = result_reg_r_22[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_68 = result_reg_r_22[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_69 = result_reg_r_22[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_70 = result_reg_r_22[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_71 = result_reg_r_22[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_72 = result_reg_r_22[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_73 = result_reg_r_22[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_74 = result_reg_r_22[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_75 = result_reg_r_22[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_76 = result_reg_r_22[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_77 = result_reg_r_22[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_78 = result_reg_r_22[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_79 = result_reg_r_22[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_80 = result_reg_r_22[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_81 = result_reg_r_22[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_82 = result_reg_r_22[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_83 = result_reg_r_22[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_84 = result_reg_r_22[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_85 = result_reg_r_22[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_86 = result_reg_r_22[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_87 = result_reg_r_22[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_88 = result_reg_r_22[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_89 = result_reg_r_22[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_90 = result_reg_r_22[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_91 = result_reg_r_22[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_92 = result_reg_r_22[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_93 = result_reg_r_22[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_94 = result_reg_r_22[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_95 = result_reg_r_22[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_96 = result_reg_r_22[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_97 = result_reg_r_22[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_98 = result_reg_r_22[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_99 = result_reg_r_22[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_100 = result_reg_r_22[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_101 = result_reg_r_22[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_102 = result_reg_r_22[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_103 = result_reg_r_22[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_104 = result_reg_r_22[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_45_105 = result_reg_r_22[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_23_hi_hi_hi_lo = {wire_res_45_98,wire_res_45_97,wire_res_45_96,wire_res_45_95,wire_res_45_94,
    wire_res_45_93,wire_res_45_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_23_hi_hi_lo_lo = {wire_res_45_84,wire_res_45_83,wire_res_45_82,wire_res_45_81,wire_res_45_80,
    wire_res_45_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_23_hi_hi_lo = {wire_res_45_91,wire_res_45_90,wire_res_45_89,wire_res_45_88,wire_res_45_87,
    wire_res_45_86,wire_res_45_85,result_reg_w_23_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_23_hi_lo_hi_lo = {wire_res_45_71,wire_res_45_70,wire_res_45_69,wire_res_45_68,wire_res_45_67,
    wire_res_45_66}; // @[BinaryDesigns2.scala 231:46]
  wire [164:0] _T_11328 = {b_aux_reg_r_22, 59'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [164:0] _GEN_1294 = {{59'd0}, a_aux_reg_r_22}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_45_59 = _GEN_1294 >= _T_11328; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_23_hi_lo_lo_lo = {wire_res_45_58,wire_res_45_57,wire_res_45_56,wire_res_45_55,wire_res_45_54,
    wire_res_45_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_23_hi_lo_lo = {wire_res_45_65,wire_res_45_64,wire_res_45_63,wire_res_45_62,wire_res_45_61,
    wire_res_45_60,wire_res_45_59,result_reg_w_23_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_23_hi_lo = {wire_res_45_78,wire_res_45_77,wire_res_45_76,wire_res_45_75,wire_res_45_74,
    wire_res_45_73,wire_res_45_72,result_reg_w_23_hi_lo_hi_lo,result_reg_w_23_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_23_hi = {wire_res_45_105,wire_res_45_104,wire_res_45_103,wire_res_45_102,wire_res_45_101,
    wire_res_45_100,wire_res_45_99,result_reg_w_23_hi_hi_hi_lo,result_reg_w_23_hi_hi_lo,result_reg_w_23_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_23_lo_hi_hi_lo = {wire_res_45_45,wire_res_45_44,wire_res_45_43,wire_res_45_42,wire_res_45_41,
    wire_res_45_40,wire_res_45_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_23_lo_hi_lo_lo = {wire_res_45_31,wire_res_45_30,wire_res_45_29,wire_res_45_28,wire_res_45_27,
    wire_res_45_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_23_lo_hi_lo = {wire_res_45_38,wire_res_45_37,wire_res_45_36,wire_res_45_35,wire_res_45_34,
    wire_res_45_33,wire_res_45_32,result_reg_w_23_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_23_lo_lo_hi_lo = {wire_res_45_18,wire_res_45_17,wire_res_45_16,wire_res_45_15,wire_res_45_14,
    wire_res_45_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_23_lo_lo_lo_lo = {wire_res_45_5,wire_res_45_4,wire_res_45_3,wire_res_45_2,wire_res_45_1,
    wire_res_45_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_23_lo_lo_lo = {wire_res_45_12,wire_res_45_11,wire_res_45_10,wire_res_45_9,wire_res_45_8,
    wire_res_45_7,wire_res_45_6,result_reg_w_23_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_23_lo_lo = {wire_res_45_25,wire_res_45_24,wire_res_45_23,wire_res_45_22,wire_res_45_21,
    wire_res_45_20,wire_res_45_19,result_reg_w_23_lo_lo_hi_lo,result_reg_w_23_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_23_lo = {wire_res_45_52,wire_res_45_51,wire_res_45_50,wire_res_45_49,wire_res_45_48,
    wire_res_45_47,wire_res_45_46,result_reg_w_23_lo_hi_hi_lo,result_reg_w_23_lo_hi_lo,result_reg_w_23_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_23 = {result_reg_w_23_hi,result_reg_w_23_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_46_0 = result_reg_w_23[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_1 = result_reg_w_23[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_2 = result_reg_w_23[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_3 = result_reg_w_23[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_4 = result_reg_w_23[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_5 = result_reg_w_23[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_6 = result_reg_w_23[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_7 = result_reg_w_23[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_8 = result_reg_w_23[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_9 = result_reg_w_23[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_10 = result_reg_w_23[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_11 = result_reg_w_23[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_12 = result_reg_w_23[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_13 = result_reg_w_23[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_14 = result_reg_w_23[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_15 = result_reg_w_23[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_16 = result_reg_w_23[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_17 = result_reg_w_23[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_18 = result_reg_w_23[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_19 = result_reg_w_23[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_20 = result_reg_w_23[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_21 = result_reg_w_23[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_22 = result_reg_w_23[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_23 = result_reg_w_23[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_24 = result_reg_w_23[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_25 = result_reg_w_23[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_26 = result_reg_w_23[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_27 = result_reg_w_23[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_28 = result_reg_w_23[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_29 = result_reg_w_23[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_30 = result_reg_w_23[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_31 = result_reg_w_23[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_32 = result_reg_w_23[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_33 = result_reg_w_23[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_34 = result_reg_w_23[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_35 = result_reg_w_23[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_36 = result_reg_w_23[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_37 = result_reg_w_23[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_38 = result_reg_w_23[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_39 = result_reg_w_23[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_40 = result_reg_w_23[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_41 = result_reg_w_23[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_42 = result_reg_w_23[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_43 = result_reg_w_23[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_44 = result_reg_w_23[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_45 = result_reg_w_23[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_46 = result_reg_w_23[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_47 = result_reg_w_23[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_48 = result_reg_w_23[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_49 = result_reg_w_23[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_50 = result_reg_w_23[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_51 = result_reg_w_23[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_52 = result_reg_w_23[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_53 = result_reg_w_23[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_54 = result_reg_w_23[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_55 = result_reg_w_23[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_56 = result_reg_w_23[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_57 = result_reg_w_23[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_59 = result_reg_w_23[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_60 = result_reg_w_23[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_61 = result_reg_w_23[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_62 = result_reg_w_23[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_63 = result_reg_w_23[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_64 = result_reg_w_23[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_65 = result_reg_w_23[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_66 = result_reg_w_23[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_67 = result_reg_w_23[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_68 = result_reg_w_23[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_69 = result_reg_w_23[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_70 = result_reg_w_23[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_71 = result_reg_w_23[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_72 = result_reg_w_23[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_73 = result_reg_w_23[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_74 = result_reg_w_23[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_75 = result_reg_w_23[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_76 = result_reg_w_23[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_77 = result_reg_w_23[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_78 = result_reg_w_23[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_79 = result_reg_w_23[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_80 = result_reg_w_23[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_81 = result_reg_w_23[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_82 = result_reg_w_23[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_83 = result_reg_w_23[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_84 = result_reg_w_23[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_85 = result_reg_w_23[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_86 = result_reg_w_23[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_87 = result_reg_w_23[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_88 = result_reg_w_23[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_89 = result_reg_w_23[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_90 = result_reg_w_23[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_91 = result_reg_w_23[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_92 = result_reg_w_23[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_93 = result_reg_w_23[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_94 = result_reg_w_23[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_95 = result_reg_w_23[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_96 = result_reg_w_23[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_97 = result_reg_w_23[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_98 = result_reg_w_23[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_99 = result_reg_w_23[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_100 = result_reg_w_23[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_101 = result_reg_w_23[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_102 = result_reg_w_23[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_103 = result_reg_w_23[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_104 = result_reg_w_23[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_46_105 = result_reg_w_23[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_0 = result_reg_r_23[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_1 = result_reg_r_23[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_2 = result_reg_r_23[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_3 = result_reg_r_23[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_4 = result_reg_r_23[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_5 = result_reg_r_23[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_6 = result_reg_r_23[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_7 = result_reg_r_23[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_8 = result_reg_r_23[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_9 = result_reg_r_23[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_10 = result_reg_r_23[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_11 = result_reg_r_23[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_12 = result_reg_r_23[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_13 = result_reg_r_23[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_14 = result_reg_r_23[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_15 = result_reg_r_23[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_16 = result_reg_r_23[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_17 = result_reg_r_23[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_18 = result_reg_r_23[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_19 = result_reg_r_23[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_20 = result_reg_r_23[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_21 = result_reg_r_23[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_22 = result_reg_r_23[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_23 = result_reg_r_23[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_24 = result_reg_r_23[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_25 = result_reg_r_23[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_26 = result_reg_r_23[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_27 = result_reg_r_23[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_28 = result_reg_r_23[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_29 = result_reg_r_23[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_30 = result_reg_r_23[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_31 = result_reg_r_23[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_32 = result_reg_r_23[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_33 = result_reg_r_23[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_34 = result_reg_r_23[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_35 = result_reg_r_23[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_36 = result_reg_r_23[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_37 = result_reg_r_23[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_38 = result_reg_r_23[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_39 = result_reg_r_23[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_40 = result_reg_r_23[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_41 = result_reg_r_23[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_42 = result_reg_r_23[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_43 = result_reg_r_23[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_44 = result_reg_r_23[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_45 = result_reg_r_23[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_46 = result_reg_r_23[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_47 = result_reg_r_23[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_48 = result_reg_r_23[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_49 = result_reg_r_23[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_50 = result_reg_r_23[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_51 = result_reg_r_23[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_52 = result_reg_r_23[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_53 = result_reg_r_23[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_54 = result_reg_r_23[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_55 = result_reg_r_23[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_56 = result_reg_r_23[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_58 = result_reg_r_23[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_59 = result_reg_r_23[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_60 = result_reg_r_23[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_61 = result_reg_r_23[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_62 = result_reg_r_23[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_63 = result_reg_r_23[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_64 = result_reg_r_23[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_65 = result_reg_r_23[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_66 = result_reg_r_23[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_67 = result_reg_r_23[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_68 = result_reg_r_23[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_69 = result_reg_r_23[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_70 = result_reg_r_23[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_71 = result_reg_r_23[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_72 = result_reg_r_23[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_73 = result_reg_r_23[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_74 = result_reg_r_23[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_75 = result_reg_r_23[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_76 = result_reg_r_23[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_77 = result_reg_r_23[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_78 = result_reg_r_23[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_79 = result_reg_r_23[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_80 = result_reg_r_23[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_81 = result_reg_r_23[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_82 = result_reg_r_23[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_83 = result_reg_r_23[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_84 = result_reg_r_23[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_85 = result_reg_r_23[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_86 = result_reg_r_23[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_87 = result_reg_r_23[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_88 = result_reg_r_23[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_89 = result_reg_r_23[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_90 = result_reg_r_23[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_91 = result_reg_r_23[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_92 = result_reg_r_23[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_93 = result_reg_r_23[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_94 = result_reg_r_23[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_95 = result_reg_r_23[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_96 = result_reg_r_23[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_97 = result_reg_r_23[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_98 = result_reg_r_23[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_99 = result_reg_r_23[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_100 = result_reg_r_23[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_101 = result_reg_r_23[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_102 = result_reg_r_23[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_103 = result_reg_r_23[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_104 = result_reg_r_23[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_47_105 = result_reg_r_23[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_24_hi_hi_hi_lo = {wire_res_47_98,wire_res_47_97,wire_res_47_96,wire_res_47_95,wire_res_47_94,
    wire_res_47_93,wire_res_47_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_24_hi_hi_lo_lo = {wire_res_47_84,wire_res_47_83,wire_res_47_82,wire_res_47_81,wire_res_47_80,
    wire_res_47_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_24_hi_hi_lo = {wire_res_47_91,wire_res_47_90,wire_res_47_89,wire_res_47_88,wire_res_47_87,
    wire_res_47_86,wire_res_47_85,result_reg_w_24_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_24_hi_lo_hi_lo = {wire_res_47_71,wire_res_47_70,wire_res_47_69,wire_res_47_68,wire_res_47_67,
    wire_res_47_66}; // @[BinaryDesigns2.scala 231:46]
  wire [162:0] _T_11332 = {b_aux_reg_r_23, 57'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [162:0] _GEN_1295 = {{57'd0}, a_aux_reg_r_23}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_47_57 = _GEN_1295 >= _T_11332; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_24_hi_lo_lo_lo = {wire_res_47_58,wire_res_47_57,wire_res_47_56,wire_res_47_55,wire_res_47_54,
    wire_res_47_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_24_hi_lo_lo = {wire_res_47_65,wire_res_47_64,wire_res_47_63,wire_res_47_62,wire_res_47_61,
    wire_res_47_60,wire_res_47_59,result_reg_w_24_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_24_hi_lo = {wire_res_47_78,wire_res_47_77,wire_res_47_76,wire_res_47_75,wire_res_47_74,
    wire_res_47_73,wire_res_47_72,result_reg_w_24_hi_lo_hi_lo,result_reg_w_24_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_24_hi = {wire_res_47_105,wire_res_47_104,wire_res_47_103,wire_res_47_102,wire_res_47_101,
    wire_res_47_100,wire_res_47_99,result_reg_w_24_hi_hi_hi_lo,result_reg_w_24_hi_hi_lo,result_reg_w_24_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_24_lo_hi_hi_lo = {wire_res_47_45,wire_res_47_44,wire_res_47_43,wire_res_47_42,wire_res_47_41,
    wire_res_47_40,wire_res_47_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_24_lo_hi_lo_lo = {wire_res_47_31,wire_res_47_30,wire_res_47_29,wire_res_47_28,wire_res_47_27,
    wire_res_47_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_24_lo_hi_lo = {wire_res_47_38,wire_res_47_37,wire_res_47_36,wire_res_47_35,wire_res_47_34,
    wire_res_47_33,wire_res_47_32,result_reg_w_24_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_24_lo_lo_hi_lo = {wire_res_47_18,wire_res_47_17,wire_res_47_16,wire_res_47_15,wire_res_47_14,
    wire_res_47_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_24_lo_lo_lo_lo = {wire_res_47_5,wire_res_47_4,wire_res_47_3,wire_res_47_2,wire_res_47_1,
    wire_res_47_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_24_lo_lo_lo = {wire_res_47_12,wire_res_47_11,wire_res_47_10,wire_res_47_9,wire_res_47_8,
    wire_res_47_7,wire_res_47_6,result_reg_w_24_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_24_lo_lo = {wire_res_47_25,wire_res_47_24,wire_res_47_23,wire_res_47_22,wire_res_47_21,
    wire_res_47_20,wire_res_47_19,result_reg_w_24_lo_lo_hi_lo,result_reg_w_24_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_24_lo = {wire_res_47_52,wire_res_47_51,wire_res_47_50,wire_res_47_49,wire_res_47_48,
    wire_res_47_47,wire_res_47_46,result_reg_w_24_lo_hi_hi_lo,result_reg_w_24_lo_hi_lo,result_reg_w_24_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_24 = {result_reg_w_24_hi,result_reg_w_24_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_48_0 = result_reg_w_24[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_1 = result_reg_w_24[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_2 = result_reg_w_24[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_3 = result_reg_w_24[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_4 = result_reg_w_24[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_5 = result_reg_w_24[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_6 = result_reg_w_24[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_7 = result_reg_w_24[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_8 = result_reg_w_24[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_9 = result_reg_w_24[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_10 = result_reg_w_24[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_11 = result_reg_w_24[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_12 = result_reg_w_24[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_13 = result_reg_w_24[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_14 = result_reg_w_24[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_15 = result_reg_w_24[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_16 = result_reg_w_24[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_17 = result_reg_w_24[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_18 = result_reg_w_24[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_19 = result_reg_w_24[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_20 = result_reg_w_24[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_21 = result_reg_w_24[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_22 = result_reg_w_24[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_23 = result_reg_w_24[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_24 = result_reg_w_24[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_25 = result_reg_w_24[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_26 = result_reg_w_24[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_27 = result_reg_w_24[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_28 = result_reg_w_24[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_29 = result_reg_w_24[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_30 = result_reg_w_24[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_31 = result_reg_w_24[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_32 = result_reg_w_24[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_33 = result_reg_w_24[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_34 = result_reg_w_24[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_35 = result_reg_w_24[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_36 = result_reg_w_24[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_37 = result_reg_w_24[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_38 = result_reg_w_24[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_39 = result_reg_w_24[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_40 = result_reg_w_24[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_41 = result_reg_w_24[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_42 = result_reg_w_24[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_43 = result_reg_w_24[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_44 = result_reg_w_24[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_45 = result_reg_w_24[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_46 = result_reg_w_24[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_47 = result_reg_w_24[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_48 = result_reg_w_24[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_49 = result_reg_w_24[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_50 = result_reg_w_24[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_51 = result_reg_w_24[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_52 = result_reg_w_24[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_53 = result_reg_w_24[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_54 = result_reg_w_24[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_55 = result_reg_w_24[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_57 = result_reg_w_24[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_58 = result_reg_w_24[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_59 = result_reg_w_24[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_60 = result_reg_w_24[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_61 = result_reg_w_24[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_62 = result_reg_w_24[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_63 = result_reg_w_24[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_64 = result_reg_w_24[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_65 = result_reg_w_24[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_66 = result_reg_w_24[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_67 = result_reg_w_24[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_68 = result_reg_w_24[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_69 = result_reg_w_24[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_70 = result_reg_w_24[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_71 = result_reg_w_24[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_72 = result_reg_w_24[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_73 = result_reg_w_24[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_74 = result_reg_w_24[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_75 = result_reg_w_24[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_76 = result_reg_w_24[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_77 = result_reg_w_24[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_78 = result_reg_w_24[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_79 = result_reg_w_24[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_80 = result_reg_w_24[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_81 = result_reg_w_24[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_82 = result_reg_w_24[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_83 = result_reg_w_24[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_84 = result_reg_w_24[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_85 = result_reg_w_24[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_86 = result_reg_w_24[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_87 = result_reg_w_24[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_88 = result_reg_w_24[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_89 = result_reg_w_24[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_90 = result_reg_w_24[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_91 = result_reg_w_24[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_92 = result_reg_w_24[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_93 = result_reg_w_24[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_94 = result_reg_w_24[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_95 = result_reg_w_24[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_96 = result_reg_w_24[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_97 = result_reg_w_24[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_98 = result_reg_w_24[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_99 = result_reg_w_24[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_100 = result_reg_w_24[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_101 = result_reg_w_24[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_102 = result_reg_w_24[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_103 = result_reg_w_24[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_104 = result_reg_w_24[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_48_105 = result_reg_w_24[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_0 = result_reg_r_24[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_1 = result_reg_r_24[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_2 = result_reg_r_24[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_3 = result_reg_r_24[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_4 = result_reg_r_24[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_5 = result_reg_r_24[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_6 = result_reg_r_24[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_7 = result_reg_r_24[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_8 = result_reg_r_24[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_9 = result_reg_r_24[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_10 = result_reg_r_24[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_11 = result_reg_r_24[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_12 = result_reg_r_24[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_13 = result_reg_r_24[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_14 = result_reg_r_24[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_15 = result_reg_r_24[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_16 = result_reg_r_24[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_17 = result_reg_r_24[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_18 = result_reg_r_24[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_19 = result_reg_r_24[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_20 = result_reg_r_24[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_21 = result_reg_r_24[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_22 = result_reg_r_24[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_23 = result_reg_r_24[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_24 = result_reg_r_24[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_25 = result_reg_r_24[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_26 = result_reg_r_24[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_27 = result_reg_r_24[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_28 = result_reg_r_24[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_29 = result_reg_r_24[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_30 = result_reg_r_24[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_31 = result_reg_r_24[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_32 = result_reg_r_24[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_33 = result_reg_r_24[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_34 = result_reg_r_24[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_35 = result_reg_r_24[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_36 = result_reg_r_24[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_37 = result_reg_r_24[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_38 = result_reg_r_24[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_39 = result_reg_r_24[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_40 = result_reg_r_24[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_41 = result_reg_r_24[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_42 = result_reg_r_24[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_43 = result_reg_r_24[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_44 = result_reg_r_24[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_45 = result_reg_r_24[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_46 = result_reg_r_24[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_47 = result_reg_r_24[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_48 = result_reg_r_24[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_49 = result_reg_r_24[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_50 = result_reg_r_24[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_51 = result_reg_r_24[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_52 = result_reg_r_24[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_53 = result_reg_r_24[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_54 = result_reg_r_24[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_56 = result_reg_r_24[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_57 = result_reg_r_24[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_58 = result_reg_r_24[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_59 = result_reg_r_24[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_60 = result_reg_r_24[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_61 = result_reg_r_24[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_62 = result_reg_r_24[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_63 = result_reg_r_24[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_64 = result_reg_r_24[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_65 = result_reg_r_24[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_66 = result_reg_r_24[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_67 = result_reg_r_24[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_68 = result_reg_r_24[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_69 = result_reg_r_24[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_70 = result_reg_r_24[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_71 = result_reg_r_24[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_72 = result_reg_r_24[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_73 = result_reg_r_24[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_74 = result_reg_r_24[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_75 = result_reg_r_24[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_76 = result_reg_r_24[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_77 = result_reg_r_24[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_78 = result_reg_r_24[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_79 = result_reg_r_24[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_80 = result_reg_r_24[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_81 = result_reg_r_24[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_82 = result_reg_r_24[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_83 = result_reg_r_24[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_84 = result_reg_r_24[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_85 = result_reg_r_24[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_86 = result_reg_r_24[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_87 = result_reg_r_24[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_88 = result_reg_r_24[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_89 = result_reg_r_24[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_90 = result_reg_r_24[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_91 = result_reg_r_24[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_92 = result_reg_r_24[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_93 = result_reg_r_24[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_94 = result_reg_r_24[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_95 = result_reg_r_24[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_96 = result_reg_r_24[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_97 = result_reg_r_24[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_98 = result_reg_r_24[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_99 = result_reg_r_24[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_100 = result_reg_r_24[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_101 = result_reg_r_24[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_102 = result_reg_r_24[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_103 = result_reg_r_24[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_104 = result_reg_r_24[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_49_105 = result_reg_r_24[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_25_hi_hi_hi_lo = {wire_res_49_98,wire_res_49_97,wire_res_49_96,wire_res_49_95,wire_res_49_94,
    wire_res_49_93,wire_res_49_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_25_hi_hi_lo_lo = {wire_res_49_84,wire_res_49_83,wire_res_49_82,wire_res_49_81,wire_res_49_80,
    wire_res_49_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_25_hi_hi_lo = {wire_res_49_91,wire_res_49_90,wire_res_49_89,wire_res_49_88,wire_res_49_87,
    wire_res_49_86,wire_res_49_85,result_reg_w_25_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_25_hi_lo_hi_lo = {wire_res_49_71,wire_res_49_70,wire_res_49_69,wire_res_49_68,wire_res_49_67,
    wire_res_49_66}; // @[BinaryDesigns2.scala 231:46]
  wire [160:0] _T_11336 = {b_aux_reg_r_24, 55'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [160:0] _GEN_1296 = {{55'd0}, a_aux_reg_r_24}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_49_55 = _GEN_1296 >= _T_11336; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_25_hi_lo_lo_lo = {wire_res_49_58,wire_res_49_57,wire_res_49_56,wire_res_49_55,wire_res_49_54,
    wire_res_49_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_25_hi_lo_lo = {wire_res_49_65,wire_res_49_64,wire_res_49_63,wire_res_49_62,wire_res_49_61,
    wire_res_49_60,wire_res_49_59,result_reg_w_25_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_25_hi_lo = {wire_res_49_78,wire_res_49_77,wire_res_49_76,wire_res_49_75,wire_res_49_74,
    wire_res_49_73,wire_res_49_72,result_reg_w_25_hi_lo_hi_lo,result_reg_w_25_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_25_hi = {wire_res_49_105,wire_res_49_104,wire_res_49_103,wire_res_49_102,wire_res_49_101,
    wire_res_49_100,wire_res_49_99,result_reg_w_25_hi_hi_hi_lo,result_reg_w_25_hi_hi_lo,result_reg_w_25_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_25_lo_hi_hi_lo = {wire_res_49_45,wire_res_49_44,wire_res_49_43,wire_res_49_42,wire_res_49_41,
    wire_res_49_40,wire_res_49_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_25_lo_hi_lo_lo = {wire_res_49_31,wire_res_49_30,wire_res_49_29,wire_res_49_28,wire_res_49_27,
    wire_res_49_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_25_lo_hi_lo = {wire_res_49_38,wire_res_49_37,wire_res_49_36,wire_res_49_35,wire_res_49_34,
    wire_res_49_33,wire_res_49_32,result_reg_w_25_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_25_lo_lo_hi_lo = {wire_res_49_18,wire_res_49_17,wire_res_49_16,wire_res_49_15,wire_res_49_14,
    wire_res_49_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_25_lo_lo_lo_lo = {wire_res_49_5,wire_res_49_4,wire_res_49_3,wire_res_49_2,wire_res_49_1,
    wire_res_49_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_25_lo_lo_lo = {wire_res_49_12,wire_res_49_11,wire_res_49_10,wire_res_49_9,wire_res_49_8,
    wire_res_49_7,wire_res_49_6,result_reg_w_25_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_25_lo_lo = {wire_res_49_25,wire_res_49_24,wire_res_49_23,wire_res_49_22,wire_res_49_21,
    wire_res_49_20,wire_res_49_19,result_reg_w_25_lo_lo_hi_lo,result_reg_w_25_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_25_lo = {wire_res_49_52,wire_res_49_51,wire_res_49_50,wire_res_49_49,wire_res_49_48,
    wire_res_49_47,wire_res_49_46,result_reg_w_25_lo_hi_hi_lo,result_reg_w_25_lo_hi_lo,result_reg_w_25_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_25 = {result_reg_w_25_hi,result_reg_w_25_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_50_0 = result_reg_w_25[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_1 = result_reg_w_25[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_2 = result_reg_w_25[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_3 = result_reg_w_25[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_4 = result_reg_w_25[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_5 = result_reg_w_25[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_6 = result_reg_w_25[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_7 = result_reg_w_25[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_8 = result_reg_w_25[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_9 = result_reg_w_25[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_10 = result_reg_w_25[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_11 = result_reg_w_25[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_12 = result_reg_w_25[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_13 = result_reg_w_25[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_14 = result_reg_w_25[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_15 = result_reg_w_25[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_16 = result_reg_w_25[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_17 = result_reg_w_25[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_18 = result_reg_w_25[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_19 = result_reg_w_25[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_20 = result_reg_w_25[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_21 = result_reg_w_25[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_22 = result_reg_w_25[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_23 = result_reg_w_25[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_24 = result_reg_w_25[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_25 = result_reg_w_25[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_26 = result_reg_w_25[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_27 = result_reg_w_25[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_28 = result_reg_w_25[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_29 = result_reg_w_25[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_30 = result_reg_w_25[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_31 = result_reg_w_25[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_32 = result_reg_w_25[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_33 = result_reg_w_25[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_34 = result_reg_w_25[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_35 = result_reg_w_25[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_36 = result_reg_w_25[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_37 = result_reg_w_25[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_38 = result_reg_w_25[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_39 = result_reg_w_25[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_40 = result_reg_w_25[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_41 = result_reg_w_25[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_42 = result_reg_w_25[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_43 = result_reg_w_25[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_44 = result_reg_w_25[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_45 = result_reg_w_25[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_46 = result_reg_w_25[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_47 = result_reg_w_25[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_48 = result_reg_w_25[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_49 = result_reg_w_25[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_50 = result_reg_w_25[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_51 = result_reg_w_25[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_52 = result_reg_w_25[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_53 = result_reg_w_25[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_55 = result_reg_w_25[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_56 = result_reg_w_25[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_57 = result_reg_w_25[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_58 = result_reg_w_25[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_59 = result_reg_w_25[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_60 = result_reg_w_25[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_61 = result_reg_w_25[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_62 = result_reg_w_25[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_63 = result_reg_w_25[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_64 = result_reg_w_25[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_65 = result_reg_w_25[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_66 = result_reg_w_25[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_67 = result_reg_w_25[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_68 = result_reg_w_25[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_69 = result_reg_w_25[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_70 = result_reg_w_25[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_71 = result_reg_w_25[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_72 = result_reg_w_25[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_73 = result_reg_w_25[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_74 = result_reg_w_25[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_75 = result_reg_w_25[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_76 = result_reg_w_25[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_77 = result_reg_w_25[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_78 = result_reg_w_25[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_79 = result_reg_w_25[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_80 = result_reg_w_25[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_81 = result_reg_w_25[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_82 = result_reg_w_25[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_83 = result_reg_w_25[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_84 = result_reg_w_25[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_85 = result_reg_w_25[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_86 = result_reg_w_25[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_87 = result_reg_w_25[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_88 = result_reg_w_25[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_89 = result_reg_w_25[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_90 = result_reg_w_25[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_91 = result_reg_w_25[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_92 = result_reg_w_25[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_93 = result_reg_w_25[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_94 = result_reg_w_25[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_95 = result_reg_w_25[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_96 = result_reg_w_25[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_97 = result_reg_w_25[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_98 = result_reg_w_25[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_99 = result_reg_w_25[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_100 = result_reg_w_25[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_101 = result_reg_w_25[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_102 = result_reg_w_25[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_103 = result_reg_w_25[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_104 = result_reg_w_25[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_50_105 = result_reg_w_25[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_0 = result_reg_r_25[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_1 = result_reg_r_25[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_2 = result_reg_r_25[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_3 = result_reg_r_25[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_4 = result_reg_r_25[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_5 = result_reg_r_25[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_6 = result_reg_r_25[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_7 = result_reg_r_25[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_8 = result_reg_r_25[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_9 = result_reg_r_25[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_10 = result_reg_r_25[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_11 = result_reg_r_25[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_12 = result_reg_r_25[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_13 = result_reg_r_25[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_14 = result_reg_r_25[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_15 = result_reg_r_25[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_16 = result_reg_r_25[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_17 = result_reg_r_25[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_18 = result_reg_r_25[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_19 = result_reg_r_25[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_20 = result_reg_r_25[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_21 = result_reg_r_25[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_22 = result_reg_r_25[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_23 = result_reg_r_25[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_24 = result_reg_r_25[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_25 = result_reg_r_25[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_26 = result_reg_r_25[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_27 = result_reg_r_25[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_28 = result_reg_r_25[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_29 = result_reg_r_25[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_30 = result_reg_r_25[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_31 = result_reg_r_25[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_32 = result_reg_r_25[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_33 = result_reg_r_25[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_34 = result_reg_r_25[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_35 = result_reg_r_25[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_36 = result_reg_r_25[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_37 = result_reg_r_25[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_38 = result_reg_r_25[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_39 = result_reg_r_25[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_40 = result_reg_r_25[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_41 = result_reg_r_25[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_42 = result_reg_r_25[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_43 = result_reg_r_25[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_44 = result_reg_r_25[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_45 = result_reg_r_25[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_46 = result_reg_r_25[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_47 = result_reg_r_25[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_48 = result_reg_r_25[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_49 = result_reg_r_25[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_50 = result_reg_r_25[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_51 = result_reg_r_25[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_52 = result_reg_r_25[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_54 = result_reg_r_25[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_55 = result_reg_r_25[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_56 = result_reg_r_25[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_57 = result_reg_r_25[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_58 = result_reg_r_25[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_59 = result_reg_r_25[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_60 = result_reg_r_25[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_61 = result_reg_r_25[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_62 = result_reg_r_25[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_63 = result_reg_r_25[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_64 = result_reg_r_25[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_65 = result_reg_r_25[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_66 = result_reg_r_25[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_67 = result_reg_r_25[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_68 = result_reg_r_25[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_69 = result_reg_r_25[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_70 = result_reg_r_25[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_71 = result_reg_r_25[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_72 = result_reg_r_25[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_73 = result_reg_r_25[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_74 = result_reg_r_25[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_75 = result_reg_r_25[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_76 = result_reg_r_25[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_77 = result_reg_r_25[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_78 = result_reg_r_25[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_79 = result_reg_r_25[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_80 = result_reg_r_25[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_81 = result_reg_r_25[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_82 = result_reg_r_25[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_83 = result_reg_r_25[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_84 = result_reg_r_25[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_85 = result_reg_r_25[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_86 = result_reg_r_25[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_87 = result_reg_r_25[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_88 = result_reg_r_25[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_89 = result_reg_r_25[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_90 = result_reg_r_25[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_91 = result_reg_r_25[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_92 = result_reg_r_25[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_93 = result_reg_r_25[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_94 = result_reg_r_25[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_95 = result_reg_r_25[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_96 = result_reg_r_25[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_97 = result_reg_r_25[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_98 = result_reg_r_25[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_99 = result_reg_r_25[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_100 = result_reg_r_25[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_101 = result_reg_r_25[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_102 = result_reg_r_25[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_103 = result_reg_r_25[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_104 = result_reg_r_25[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_51_105 = result_reg_r_25[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_26_hi_hi_hi_lo = {wire_res_51_98,wire_res_51_97,wire_res_51_96,wire_res_51_95,wire_res_51_94,
    wire_res_51_93,wire_res_51_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_26_hi_hi_lo_lo = {wire_res_51_84,wire_res_51_83,wire_res_51_82,wire_res_51_81,wire_res_51_80,
    wire_res_51_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_26_hi_hi_lo = {wire_res_51_91,wire_res_51_90,wire_res_51_89,wire_res_51_88,wire_res_51_87,
    wire_res_51_86,wire_res_51_85,result_reg_w_26_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_26_hi_lo_hi_lo = {wire_res_51_71,wire_res_51_70,wire_res_51_69,wire_res_51_68,wire_res_51_67,
    wire_res_51_66}; // @[BinaryDesigns2.scala 231:46]
  wire [158:0] _T_11340 = {b_aux_reg_r_25, 53'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [158:0] _GEN_1297 = {{53'd0}, a_aux_reg_r_25}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_51_53 = _GEN_1297 >= _T_11340; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_26_hi_lo_lo_lo = {wire_res_51_58,wire_res_51_57,wire_res_51_56,wire_res_51_55,wire_res_51_54,
    wire_res_51_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_26_hi_lo_lo = {wire_res_51_65,wire_res_51_64,wire_res_51_63,wire_res_51_62,wire_res_51_61,
    wire_res_51_60,wire_res_51_59,result_reg_w_26_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_26_hi_lo = {wire_res_51_78,wire_res_51_77,wire_res_51_76,wire_res_51_75,wire_res_51_74,
    wire_res_51_73,wire_res_51_72,result_reg_w_26_hi_lo_hi_lo,result_reg_w_26_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_26_hi = {wire_res_51_105,wire_res_51_104,wire_res_51_103,wire_res_51_102,wire_res_51_101,
    wire_res_51_100,wire_res_51_99,result_reg_w_26_hi_hi_hi_lo,result_reg_w_26_hi_hi_lo,result_reg_w_26_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_26_lo_hi_hi_lo = {wire_res_51_45,wire_res_51_44,wire_res_51_43,wire_res_51_42,wire_res_51_41,
    wire_res_51_40,wire_res_51_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_26_lo_hi_lo_lo = {wire_res_51_31,wire_res_51_30,wire_res_51_29,wire_res_51_28,wire_res_51_27,
    wire_res_51_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_26_lo_hi_lo = {wire_res_51_38,wire_res_51_37,wire_res_51_36,wire_res_51_35,wire_res_51_34,
    wire_res_51_33,wire_res_51_32,result_reg_w_26_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_26_lo_lo_hi_lo = {wire_res_51_18,wire_res_51_17,wire_res_51_16,wire_res_51_15,wire_res_51_14,
    wire_res_51_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_26_lo_lo_lo_lo = {wire_res_51_5,wire_res_51_4,wire_res_51_3,wire_res_51_2,wire_res_51_1,
    wire_res_51_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_26_lo_lo_lo = {wire_res_51_12,wire_res_51_11,wire_res_51_10,wire_res_51_9,wire_res_51_8,
    wire_res_51_7,wire_res_51_6,result_reg_w_26_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_26_lo_lo = {wire_res_51_25,wire_res_51_24,wire_res_51_23,wire_res_51_22,wire_res_51_21,
    wire_res_51_20,wire_res_51_19,result_reg_w_26_lo_lo_hi_lo,result_reg_w_26_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_26_lo = {wire_res_51_52,wire_res_51_51,wire_res_51_50,wire_res_51_49,wire_res_51_48,
    wire_res_51_47,wire_res_51_46,result_reg_w_26_lo_hi_hi_lo,result_reg_w_26_lo_hi_lo,result_reg_w_26_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_26 = {result_reg_w_26_hi,result_reg_w_26_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_52_0 = result_reg_w_26[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_1 = result_reg_w_26[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_2 = result_reg_w_26[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_3 = result_reg_w_26[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_4 = result_reg_w_26[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_5 = result_reg_w_26[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_6 = result_reg_w_26[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_7 = result_reg_w_26[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_8 = result_reg_w_26[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_9 = result_reg_w_26[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_10 = result_reg_w_26[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_11 = result_reg_w_26[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_12 = result_reg_w_26[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_13 = result_reg_w_26[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_14 = result_reg_w_26[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_15 = result_reg_w_26[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_16 = result_reg_w_26[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_17 = result_reg_w_26[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_18 = result_reg_w_26[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_19 = result_reg_w_26[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_20 = result_reg_w_26[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_21 = result_reg_w_26[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_22 = result_reg_w_26[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_23 = result_reg_w_26[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_24 = result_reg_w_26[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_25 = result_reg_w_26[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_26 = result_reg_w_26[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_27 = result_reg_w_26[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_28 = result_reg_w_26[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_29 = result_reg_w_26[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_30 = result_reg_w_26[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_31 = result_reg_w_26[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_32 = result_reg_w_26[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_33 = result_reg_w_26[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_34 = result_reg_w_26[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_35 = result_reg_w_26[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_36 = result_reg_w_26[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_37 = result_reg_w_26[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_38 = result_reg_w_26[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_39 = result_reg_w_26[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_40 = result_reg_w_26[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_41 = result_reg_w_26[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_42 = result_reg_w_26[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_43 = result_reg_w_26[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_44 = result_reg_w_26[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_45 = result_reg_w_26[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_46 = result_reg_w_26[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_47 = result_reg_w_26[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_48 = result_reg_w_26[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_49 = result_reg_w_26[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_50 = result_reg_w_26[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_51 = result_reg_w_26[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_53 = result_reg_w_26[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_54 = result_reg_w_26[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_55 = result_reg_w_26[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_56 = result_reg_w_26[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_57 = result_reg_w_26[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_58 = result_reg_w_26[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_59 = result_reg_w_26[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_60 = result_reg_w_26[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_61 = result_reg_w_26[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_62 = result_reg_w_26[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_63 = result_reg_w_26[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_64 = result_reg_w_26[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_65 = result_reg_w_26[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_66 = result_reg_w_26[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_67 = result_reg_w_26[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_68 = result_reg_w_26[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_69 = result_reg_w_26[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_70 = result_reg_w_26[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_71 = result_reg_w_26[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_72 = result_reg_w_26[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_73 = result_reg_w_26[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_74 = result_reg_w_26[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_75 = result_reg_w_26[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_76 = result_reg_w_26[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_77 = result_reg_w_26[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_78 = result_reg_w_26[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_79 = result_reg_w_26[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_80 = result_reg_w_26[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_81 = result_reg_w_26[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_82 = result_reg_w_26[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_83 = result_reg_w_26[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_84 = result_reg_w_26[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_85 = result_reg_w_26[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_86 = result_reg_w_26[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_87 = result_reg_w_26[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_88 = result_reg_w_26[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_89 = result_reg_w_26[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_90 = result_reg_w_26[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_91 = result_reg_w_26[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_92 = result_reg_w_26[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_93 = result_reg_w_26[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_94 = result_reg_w_26[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_95 = result_reg_w_26[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_96 = result_reg_w_26[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_97 = result_reg_w_26[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_98 = result_reg_w_26[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_99 = result_reg_w_26[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_100 = result_reg_w_26[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_101 = result_reg_w_26[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_102 = result_reg_w_26[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_103 = result_reg_w_26[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_104 = result_reg_w_26[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_52_105 = result_reg_w_26[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_0 = result_reg_r_26[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_1 = result_reg_r_26[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_2 = result_reg_r_26[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_3 = result_reg_r_26[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_4 = result_reg_r_26[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_5 = result_reg_r_26[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_6 = result_reg_r_26[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_7 = result_reg_r_26[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_8 = result_reg_r_26[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_9 = result_reg_r_26[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_10 = result_reg_r_26[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_11 = result_reg_r_26[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_12 = result_reg_r_26[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_13 = result_reg_r_26[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_14 = result_reg_r_26[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_15 = result_reg_r_26[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_16 = result_reg_r_26[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_17 = result_reg_r_26[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_18 = result_reg_r_26[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_19 = result_reg_r_26[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_20 = result_reg_r_26[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_21 = result_reg_r_26[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_22 = result_reg_r_26[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_23 = result_reg_r_26[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_24 = result_reg_r_26[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_25 = result_reg_r_26[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_26 = result_reg_r_26[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_27 = result_reg_r_26[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_28 = result_reg_r_26[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_29 = result_reg_r_26[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_30 = result_reg_r_26[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_31 = result_reg_r_26[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_32 = result_reg_r_26[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_33 = result_reg_r_26[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_34 = result_reg_r_26[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_35 = result_reg_r_26[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_36 = result_reg_r_26[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_37 = result_reg_r_26[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_38 = result_reg_r_26[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_39 = result_reg_r_26[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_40 = result_reg_r_26[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_41 = result_reg_r_26[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_42 = result_reg_r_26[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_43 = result_reg_r_26[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_44 = result_reg_r_26[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_45 = result_reg_r_26[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_46 = result_reg_r_26[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_47 = result_reg_r_26[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_48 = result_reg_r_26[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_49 = result_reg_r_26[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_50 = result_reg_r_26[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_52 = result_reg_r_26[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_53 = result_reg_r_26[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_54 = result_reg_r_26[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_55 = result_reg_r_26[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_56 = result_reg_r_26[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_57 = result_reg_r_26[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_58 = result_reg_r_26[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_59 = result_reg_r_26[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_60 = result_reg_r_26[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_61 = result_reg_r_26[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_62 = result_reg_r_26[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_63 = result_reg_r_26[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_64 = result_reg_r_26[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_65 = result_reg_r_26[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_66 = result_reg_r_26[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_67 = result_reg_r_26[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_68 = result_reg_r_26[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_69 = result_reg_r_26[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_70 = result_reg_r_26[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_71 = result_reg_r_26[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_72 = result_reg_r_26[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_73 = result_reg_r_26[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_74 = result_reg_r_26[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_75 = result_reg_r_26[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_76 = result_reg_r_26[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_77 = result_reg_r_26[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_78 = result_reg_r_26[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_79 = result_reg_r_26[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_80 = result_reg_r_26[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_81 = result_reg_r_26[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_82 = result_reg_r_26[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_83 = result_reg_r_26[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_84 = result_reg_r_26[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_85 = result_reg_r_26[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_86 = result_reg_r_26[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_87 = result_reg_r_26[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_88 = result_reg_r_26[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_89 = result_reg_r_26[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_90 = result_reg_r_26[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_91 = result_reg_r_26[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_92 = result_reg_r_26[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_93 = result_reg_r_26[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_94 = result_reg_r_26[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_95 = result_reg_r_26[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_96 = result_reg_r_26[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_97 = result_reg_r_26[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_98 = result_reg_r_26[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_99 = result_reg_r_26[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_100 = result_reg_r_26[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_101 = result_reg_r_26[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_102 = result_reg_r_26[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_103 = result_reg_r_26[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_104 = result_reg_r_26[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_53_105 = result_reg_r_26[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_27_hi_hi_hi_lo = {wire_res_53_98,wire_res_53_97,wire_res_53_96,wire_res_53_95,wire_res_53_94,
    wire_res_53_93,wire_res_53_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_27_hi_hi_lo_lo = {wire_res_53_84,wire_res_53_83,wire_res_53_82,wire_res_53_81,wire_res_53_80,
    wire_res_53_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_27_hi_hi_lo = {wire_res_53_91,wire_res_53_90,wire_res_53_89,wire_res_53_88,wire_res_53_87,
    wire_res_53_86,wire_res_53_85,result_reg_w_27_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_27_hi_lo_hi_lo = {wire_res_53_71,wire_res_53_70,wire_res_53_69,wire_res_53_68,wire_res_53_67,
    wire_res_53_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_27_hi_lo_lo_lo = {wire_res_53_58,wire_res_53_57,wire_res_53_56,wire_res_53_55,wire_res_53_54,
    wire_res_53_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_27_hi_lo_lo = {wire_res_53_65,wire_res_53_64,wire_res_53_63,wire_res_53_62,wire_res_53_61,
    wire_res_53_60,wire_res_53_59,result_reg_w_27_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_27_hi_lo = {wire_res_53_78,wire_res_53_77,wire_res_53_76,wire_res_53_75,wire_res_53_74,
    wire_res_53_73,wire_res_53_72,result_reg_w_27_hi_lo_hi_lo,result_reg_w_27_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_27_hi = {wire_res_53_105,wire_res_53_104,wire_res_53_103,wire_res_53_102,wire_res_53_101,
    wire_res_53_100,wire_res_53_99,result_reg_w_27_hi_hi_hi_lo,result_reg_w_27_hi_hi_lo,result_reg_w_27_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [156:0] _T_11344 = {b_aux_reg_r_26, 51'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [156:0] _GEN_1298 = {{51'd0}, a_aux_reg_r_26}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_53_51 = _GEN_1298 >= _T_11344; // @[BinaryDesigns2.scala 224:35]
  wire [6:0] result_reg_w_27_lo_hi_hi_lo = {wire_res_53_45,wire_res_53_44,wire_res_53_43,wire_res_53_42,wire_res_53_41,
    wire_res_53_40,wire_res_53_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_27_lo_hi_lo_lo = {wire_res_53_31,wire_res_53_30,wire_res_53_29,wire_res_53_28,wire_res_53_27,
    wire_res_53_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_27_lo_hi_lo = {wire_res_53_38,wire_res_53_37,wire_res_53_36,wire_res_53_35,wire_res_53_34,
    wire_res_53_33,wire_res_53_32,result_reg_w_27_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_27_lo_lo_hi_lo = {wire_res_53_18,wire_res_53_17,wire_res_53_16,wire_res_53_15,wire_res_53_14,
    wire_res_53_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_27_lo_lo_lo_lo = {wire_res_53_5,wire_res_53_4,wire_res_53_3,wire_res_53_2,wire_res_53_1,
    wire_res_53_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_27_lo_lo_lo = {wire_res_53_12,wire_res_53_11,wire_res_53_10,wire_res_53_9,wire_res_53_8,
    wire_res_53_7,wire_res_53_6,result_reg_w_27_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_27_lo_lo = {wire_res_53_25,wire_res_53_24,wire_res_53_23,wire_res_53_22,wire_res_53_21,
    wire_res_53_20,wire_res_53_19,result_reg_w_27_lo_lo_hi_lo,result_reg_w_27_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_27_lo = {wire_res_53_52,wire_res_53_51,wire_res_53_50,wire_res_53_49,wire_res_53_48,
    wire_res_53_47,wire_res_53_46,result_reg_w_27_lo_hi_hi_lo,result_reg_w_27_lo_hi_lo,result_reg_w_27_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_27 = {result_reg_w_27_hi,result_reg_w_27_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_54_0 = result_reg_w_27[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_1 = result_reg_w_27[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_2 = result_reg_w_27[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_3 = result_reg_w_27[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_4 = result_reg_w_27[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_5 = result_reg_w_27[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_6 = result_reg_w_27[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_7 = result_reg_w_27[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_8 = result_reg_w_27[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_9 = result_reg_w_27[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_10 = result_reg_w_27[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_11 = result_reg_w_27[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_12 = result_reg_w_27[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_13 = result_reg_w_27[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_14 = result_reg_w_27[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_15 = result_reg_w_27[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_16 = result_reg_w_27[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_17 = result_reg_w_27[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_18 = result_reg_w_27[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_19 = result_reg_w_27[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_20 = result_reg_w_27[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_21 = result_reg_w_27[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_22 = result_reg_w_27[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_23 = result_reg_w_27[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_24 = result_reg_w_27[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_25 = result_reg_w_27[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_26 = result_reg_w_27[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_27 = result_reg_w_27[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_28 = result_reg_w_27[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_29 = result_reg_w_27[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_30 = result_reg_w_27[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_31 = result_reg_w_27[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_32 = result_reg_w_27[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_33 = result_reg_w_27[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_34 = result_reg_w_27[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_35 = result_reg_w_27[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_36 = result_reg_w_27[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_37 = result_reg_w_27[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_38 = result_reg_w_27[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_39 = result_reg_w_27[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_40 = result_reg_w_27[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_41 = result_reg_w_27[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_42 = result_reg_w_27[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_43 = result_reg_w_27[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_44 = result_reg_w_27[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_45 = result_reg_w_27[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_46 = result_reg_w_27[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_47 = result_reg_w_27[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_48 = result_reg_w_27[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_49 = result_reg_w_27[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_51 = result_reg_w_27[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_52 = result_reg_w_27[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_53 = result_reg_w_27[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_54 = result_reg_w_27[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_55 = result_reg_w_27[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_56 = result_reg_w_27[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_57 = result_reg_w_27[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_58 = result_reg_w_27[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_59 = result_reg_w_27[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_60 = result_reg_w_27[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_61 = result_reg_w_27[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_62 = result_reg_w_27[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_63 = result_reg_w_27[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_64 = result_reg_w_27[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_65 = result_reg_w_27[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_66 = result_reg_w_27[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_67 = result_reg_w_27[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_68 = result_reg_w_27[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_69 = result_reg_w_27[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_70 = result_reg_w_27[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_71 = result_reg_w_27[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_72 = result_reg_w_27[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_73 = result_reg_w_27[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_74 = result_reg_w_27[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_75 = result_reg_w_27[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_76 = result_reg_w_27[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_77 = result_reg_w_27[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_78 = result_reg_w_27[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_79 = result_reg_w_27[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_80 = result_reg_w_27[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_81 = result_reg_w_27[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_82 = result_reg_w_27[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_83 = result_reg_w_27[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_84 = result_reg_w_27[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_85 = result_reg_w_27[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_86 = result_reg_w_27[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_87 = result_reg_w_27[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_88 = result_reg_w_27[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_89 = result_reg_w_27[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_90 = result_reg_w_27[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_91 = result_reg_w_27[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_92 = result_reg_w_27[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_93 = result_reg_w_27[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_94 = result_reg_w_27[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_95 = result_reg_w_27[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_96 = result_reg_w_27[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_97 = result_reg_w_27[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_98 = result_reg_w_27[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_99 = result_reg_w_27[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_100 = result_reg_w_27[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_101 = result_reg_w_27[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_102 = result_reg_w_27[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_103 = result_reg_w_27[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_104 = result_reg_w_27[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_54_105 = result_reg_w_27[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_0 = result_reg_r_27[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_1 = result_reg_r_27[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_2 = result_reg_r_27[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_3 = result_reg_r_27[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_4 = result_reg_r_27[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_5 = result_reg_r_27[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_6 = result_reg_r_27[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_7 = result_reg_r_27[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_8 = result_reg_r_27[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_9 = result_reg_r_27[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_10 = result_reg_r_27[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_11 = result_reg_r_27[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_12 = result_reg_r_27[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_13 = result_reg_r_27[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_14 = result_reg_r_27[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_15 = result_reg_r_27[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_16 = result_reg_r_27[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_17 = result_reg_r_27[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_18 = result_reg_r_27[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_19 = result_reg_r_27[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_20 = result_reg_r_27[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_21 = result_reg_r_27[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_22 = result_reg_r_27[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_23 = result_reg_r_27[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_24 = result_reg_r_27[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_25 = result_reg_r_27[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_26 = result_reg_r_27[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_27 = result_reg_r_27[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_28 = result_reg_r_27[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_29 = result_reg_r_27[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_30 = result_reg_r_27[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_31 = result_reg_r_27[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_32 = result_reg_r_27[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_33 = result_reg_r_27[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_34 = result_reg_r_27[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_35 = result_reg_r_27[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_36 = result_reg_r_27[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_37 = result_reg_r_27[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_38 = result_reg_r_27[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_39 = result_reg_r_27[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_40 = result_reg_r_27[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_41 = result_reg_r_27[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_42 = result_reg_r_27[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_43 = result_reg_r_27[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_44 = result_reg_r_27[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_45 = result_reg_r_27[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_46 = result_reg_r_27[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_47 = result_reg_r_27[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_48 = result_reg_r_27[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_50 = result_reg_r_27[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_51 = result_reg_r_27[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_52 = result_reg_r_27[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_53 = result_reg_r_27[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_54 = result_reg_r_27[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_55 = result_reg_r_27[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_56 = result_reg_r_27[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_57 = result_reg_r_27[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_58 = result_reg_r_27[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_59 = result_reg_r_27[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_60 = result_reg_r_27[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_61 = result_reg_r_27[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_62 = result_reg_r_27[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_63 = result_reg_r_27[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_64 = result_reg_r_27[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_65 = result_reg_r_27[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_66 = result_reg_r_27[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_67 = result_reg_r_27[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_68 = result_reg_r_27[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_69 = result_reg_r_27[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_70 = result_reg_r_27[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_71 = result_reg_r_27[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_72 = result_reg_r_27[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_73 = result_reg_r_27[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_74 = result_reg_r_27[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_75 = result_reg_r_27[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_76 = result_reg_r_27[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_77 = result_reg_r_27[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_78 = result_reg_r_27[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_79 = result_reg_r_27[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_80 = result_reg_r_27[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_81 = result_reg_r_27[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_82 = result_reg_r_27[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_83 = result_reg_r_27[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_84 = result_reg_r_27[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_85 = result_reg_r_27[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_86 = result_reg_r_27[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_87 = result_reg_r_27[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_88 = result_reg_r_27[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_89 = result_reg_r_27[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_90 = result_reg_r_27[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_91 = result_reg_r_27[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_92 = result_reg_r_27[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_93 = result_reg_r_27[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_94 = result_reg_r_27[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_95 = result_reg_r_27[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_96 = result_reg_r_27[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_97 = result_reg_r_27[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_98 = result_reg_r_27[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_99 = result_reg_r_27[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_100 = result_reg_r_27[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_101 = result_reg_r_27[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_102 = result_reg_r_27[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_103 = result_reg_r_27[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_104 = result_reg_r_27[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_55_105 = result_reg_r_27[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_28_hi_hi_hi_lo = {wire_res_55_98,wire_res_55_97,wire_res_55_96,wire_res_55_95,wire_res_55_94,
    wire_res_55_93,wire_res_55_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_28_hi_hi_lo_lo = {wire_res_55_84,wire_res_55_83,wire_res_55_82,wire_res_55_81,wire_res_55_80,
    wire_res_55_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_28_hi_hi_lo = {wire_res_55_91,wire_res_55_90,wire_res_55_89,wire_res_55_88,wire_res_55_87,
    wire_res_55_86,wire_res_55_85,result_reg_w_28_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_28_hi_lo_hi_lo = {wire_res_55_71,wire_res_55_70,wire_res_55_69,wire_res_55_68,wire_res_55_67,
    wire_res_55_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_28_hi_lo_lo_lo = {wire_res_55_58,wire_res_55_57,wire_res_55_56,wire_res_55_55,wire_res_55_54,
    wire_res_55_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_28_hi_lo_lo = {wire_res_55_65,wire_res_55_64,wire_res_55_63,wire_res_55_62,wire_res_55_61,
    wire_res_55_60,wire_res_55_59,result_reg_w_28_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_28_hi_lo = {wire_res_55_78,wire_res_55_77,wire_res_55_76,wire_res_55_75,wire_res_55_74,
    wire_res_55_73,wire_res_55_72,result_reg_w_28_hi_lo_hi_lo,result_reg_w_28_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_28_hi = {wire_res_55_105,wire_res_55_104,wire_res_55_103,wire_res_55_102,wire_res_55_101,
    wire_res_55_100,wire_res_55_99,result_reg_w_28_hi_hi_hi_lo,result_reg_w_28_hi_hi_lo,result_reg_w_28_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [154:0] _T_11348 = {b_aux_reg_r_27, 49'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [154:0] _GEN_1299 = {{49'd0}, a_aux_reg_r_27}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_55_49 = _GEN_1299 >= _T_11348; // @[BinaryDesigns2.scala 224:35]
  wire [6:0] result_reg_w_28_lo_hi_hi_lo = {wire_res_55_45,wire_res_55_44,wire_res_55_43,wire_res_55_42,wire_res_55_41,
    wire_res_55_40,wire_res_55_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_28_lo_hi_lo_lo = {wire_res_55_31,wire_res_55_30,wire_res_55_29,wire_res_55_28,wire_res_55_27,
    wire_res_55_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_28_lo_hi_lo = {wire_res_55_38,wire_res_55_37,wire_res_55_36,wire_res_55_35,wire_res_55_34,
    wire_res_55_33,wire_res_55_32,result_reg_w_28_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_28_lo_lo_hi_lo = {wire_res_55_18,wire_res_55_17,wire_res_55_16,wire_res_55_15,wire_res_55_14,
    wire_res_55_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_28_lo_lo_lo_lo = {wire_res_55_5,wire_res_55_4,wire_res_55_3,wire_res_55_2,wire_res_55_1,
    wire_res_55_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_28_lo_lo_lo = {wire_res_55_12,wire_res_55_11,wire_res_55_10,wire_res_55_9,wire_res_55_8,
    wire_res_55_7,wire_res_55_6,result_reg_w_28_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_28_lo_lo = {wire_res_55_25,wire_res_55_24,wire_res_55_23,wire_res_55_22,wire_res_55_21,
    wire_res_55_20,wire_res_55_19,result_reg_w_28_lo_lo_hi_lo,result_reg_w_28_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_28_lo = {wire_res_55_52,wire_res_55_51,wire_res_55_50,wire_res_55_49,wire_res_55_48,
    wire_res_55_47,wire_res_55_46,result_reg_w_28_lo_hi_hi_lo,result_reg_w_28_lo_hi_lo,result_reg_w_28_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_28 = {result_reg_w_28_hi,result_reg_w_28_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_56_0 = result_reg_w_28[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_1 = result_reg_w_28[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_2 = result_reg_w_28[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_3 = result_reg_w_28[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_4 = result_reg_w_28[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_5 = result_reg_w_28[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_6 = result_reg_w_28[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_7 = result_reg_w_28[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_8 = result_reg_w_28[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_9 = result_reg_w_28[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_10 = result_reg_w_28[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_11 = result_reg_w_28[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_12 = result_reg_w_28[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_13 = result_reg_w_28[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_14 = result_reg_w_28[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_15 = result_reg_w_28[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_16 = result_reg_w_28[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_17 = result_reg_w_28[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_18 = result_reg_w_28[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_19 = result_reg_w_28[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_20 = result_reg_w_28[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_21 = result_reg_w_28[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_22 = result_reg_w_28[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_23 = result_reg_w_28[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_24 = result_reg_w_28[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_25 = result_reg_w_28[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_26 = result_reg_w_28[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_27 = result_reg_w_28[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_28 = result_reg_w_28[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_29 = result_reg_w_28[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_30 = result_reg_w_28[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_31 = result_reg_w_28[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_32 = result_reg_w_28[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_33 = result_reg_w_28[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_34 = result_reg_w_28[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_35 = result_reg_w_28[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_36 = result_reg_w_28[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_37 = result_reg_w_28[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_38 = result_reg_w_28[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_39 = result_reg_w_28[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_40 = result_reg_w_28[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_41 = result_reg_w_28[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_42 = result_reg_w_28[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_43 = result_reg_w_28[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_44 = result_reg_w_28[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_45 = result_reg_w_28[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_46 = result_reg_w_28[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_47 = result_reg_w_28[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_49 = result_reg_w_28[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_50 = result_reg_w_28[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_51 = result_reg_w_28[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_52 = result_reg_w_28[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_53 = result_reg_w_28[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_54 = result_reg_w_28[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_55 = result_reg_w_28[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_56 = result_reg_w_28[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_57 = result_reg_w_28[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_58 = result_reg_w_28[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_59 = result_reg_w_28[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_60 = result_reg_w_28[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_61 = result_reg_w_28[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_62 = result_reg_w_28[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_63 = result_reg_w_28[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_64 = result_reg_w_28[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_65 = result_reg_w_28[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_66 = result_reg_w_28[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_67 = result_reg_w_28[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_68 = result_reg_w_28[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_69 = result_reg_w_28[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_70 = result_reg_w_28[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_71 = result_reg_w_28[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_72 = result_reg_w_28[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_73 = result_reg_w_28[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_74 = result_reg_w_28[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_75 = result_reg_w_28[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_76 = result_reg_w_28[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_77 = result_reg_w_28[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_78 = result_reg_w_28[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_79 = result_reg_w_28[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_80 = result_reg_w_28[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_81 = result_reg_w_28[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_82 = result_reg_w_28[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_83 = result_reg_w_28[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_84 = result_reg_w_28[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_85 = result_reg_w_28[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_86 = result_reg_w_28[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_87 = result_reg_w_28[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_88 = result_reg_w_28[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_89 = result_reg_w_28[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_90 = result_reg_w_28[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_91 = result_reg_w_28[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_92 = result_reg_w_28[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_93 = result_reg_w_28[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_94 = result_reg_w_28[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_95 = result_reg_w_28[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_96 = result_reg_w_28[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_97 = result_reg_w_28[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_98 = result_reg_w_28[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_99 = result_reg_w_28[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_100 = result_reg_w_28[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_101 = result_reg_w_28[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_102 = result_reg_w_28[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_103 = result_reg_w_28[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_104 = result_reg_w_28[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_56_105 = result_reg_w_28[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_0 = result_reg_r_28[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_1 = result_reg_r_28[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_2 = result_reg_r_28[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_3 = result_reg_r_28[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_4 = result_reg_r_28[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_5 = result_reg_r_28[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_6 = result_reg_r_28[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_7 = result_reg_r_28[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_8 = result_reg_r_28[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_9 = result_reg_r_28[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_10 = result_reg_r_28[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_11 = result_reg_r_28[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_12 = result_reg_r_28[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_13 = result_reg_r_28[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_14 = result_reg_r_28[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_15 = result_reg_r_28[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_16 = result_reg_r_28[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_17 = result_reg_r_28[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_18 = result_reg_r_28[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_19 = result_reg_r_28[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_20 = result_reg_r_28[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_21 = result_reg_r_28[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_22 = result_reg_r_28[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_23 = result_reg_r_28[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_24 = result_reg_r_28[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_25 = result_reg_r_28[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_26 = result_reg_r_28[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_27 = result_reg_r_28[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_28 = result_reg_r_28[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_29 = result_reg_r_28[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_30 = result_reg_r_28[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_31 = result_reg_r_28[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_32 = result_reg_r_28[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_33 = result_reg_r_28[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_34 = result_reg_r_28[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_35 = result_reg_r_28[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_36 = result_reg_r_28[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_37 = result_reg_r_28[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_38 = result_reg_r_28[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_39 = result_reg_r_28[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_40 = result_reg_r_28[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_41 = result_reg_r_28[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_42 = result_reg_r_28[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_43 = result_reg_r_28[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_44 = result_reg_r_28[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_45 = result_reg_r_28[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_46 = result_reg_r_28[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_48 = result_reg_r_28[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_49 = result_reg_r_28[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_50 = result_reg_r_28[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_51 = result_reg_r_28[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_52 = result_reg_r_28[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_53 = result_reg_r_28[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_54 = result_reg_r_28[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_55 = result_reg_r_28[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_56 = result_reg_r_28[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_57 = result_reg_r_28[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_58 = result_reg_r_28[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_59 = result_reg_r_28[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_60 = result_reg_r_28[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_61 = result_reg_r_28[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_62 = result_reg_r_28[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_63 = result_reg_r_28[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_64 = result_reg_r_28[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_65 = result_reg_r_28[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_66 = result_reg_r_28[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_67 = result_reg_r_28[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_68 = result_reg_r_28[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_69 = result_reg_r_28[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_70 = result_reg_r_28[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_71 = result_reg_r_28[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_72 = result_reg_r_28[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_73 = result_reg_r_28[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_74 = result_reg_r_28[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_75 = result_reg_r_28[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_76 = result_reg_r_28[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_77 = result_reg_r_28[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_78 = result_reg_r_28[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_79 = result_reg_r_28[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_80 = result_reg_r_28[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_81 = result_reg_r_28[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_82 = result_reg_r_28[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_83 = result_reg_r_28[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_84 = result_reg_r_28[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_85 = result_reg_r_28[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_86 = result_reg_r_28[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_87 = result_reg_r_28[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_88 = result_reg_r_28[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_89 = result_reg_r_28[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_90 = result_reg_r_28[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_91 = result_reg_r_28[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_92 = result_reg_r_28[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_93 = result_reg_r_28[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_94 = result_reg_r_28[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_95 = result_reg_r_28[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_96 = result_reg_r_28[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_97 = result_reg_r_28[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_98 = result_reg_r_28[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_99 = result_reg_r_28[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_100 = result_reg_r_28[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_101 = result_reg_r_28[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_102 = result_reg_r_28[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_103 = result_reg_r_28[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_104 = result_reg_r_28[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_57_105 = result_reg_r_28[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_29_hi_hi_hi_lo = {wire_res_57_98,wire_res_57_97,wire_res_57_96,wire_res_57_95,wire_res_57_94,
    wire_res_57_93,wire_res_57_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_29_hi_hi_lo_lo = {wire_res_57_84,wire_res_57_83,wire_res_57_82,wire_res_57_81,wire_res_57_80,
    wire_res_57_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_29_hi_hi_lo = {wire_res_57_91,wire_res_57_90,wire_res_57_89,wire_res_57_88,wire_res_57_87,
    wire_res_57_86,wire_res_57_85,result_reg_w_29_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_29_hi_lo_hi_lo = {wire_res_57_71,wire_res_57_70,wire_res_57_69,wire_res_57_68,wire_res_57_67,
    wire_res_57_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_29_hi_lo_lo_lo = {wire_res_57_58,wire_res_57_57,wire_res_57_56,wire_res_57_55,wire_res_57_54,
    wire_res_57_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_29_hi_lo_lo = {wire_res_57_65,wire_res_57_64,wire_res_57_63,wire_res_57_62,wire_res_57_61,
    wire_res_57_60,wire_res_57_59,result_reg_w_29_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_29_hi_lo = {wire_res_57_78,wire_res_57_77,wire_res_57_76,wire_res_57_75,wire_res_57_74,
    wire_res_57_73,wire_res_57_72,result_reg_w_29_hi_lo_hi_lo,result_reg_w_29_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_29_hi = {wire_res_57_105,wire_res_57_104,wire_res_57_103,wire_res_57_102,wire_res_57_101,
    wire_res_57_100,wire_res_57_99,result_reg_w_29_hi_hi_hi_lo,result_reg_w_29_hi_hi_lo,result_reg_w_29_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [152:0] _T_11352 = {b_aux_reg_r_28, 47'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [152:0] _GEN_1300 = {{47'd0}, a_aux_reg_r_28}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_57_47 = _GEN_1300 >= _T_11352; // @[BinaryDesigns2.scala 224:35]
  wire [6:0] result_reg_w_29_lo_hi_hi_lo = {wire_res_57_45,wire_res_57_44,wire_res_57_43,wire_res_57_42,wire_res_57_41,
    wire_res_57_40,wire_res_57_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_29_lo_hi_lo_lo = {wire_res_57_31,wire_res_57_30,wire_res_57_29,wire_res_57_28,wire_res_57_27,
    wire_res_57_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_29_lo_hi_lo = {wire_res_57_38,wire_res_57_37,wire_res_57_36,wire_res_57_35,wire_res_57_34,
    wire_res_57_33,wire_res_57_32,result_reg_w_29_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_29_lo_lo_hi_lo = {wire_res_57_18,wire_res_57_17,wire_res_57_16,wire_res_57_15,wire_res_57_14,
    wire_res_57_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_29_lo_lo_lo_lo = {wire_res_57_5,wire_res_57_4,wire_res_57_3,wire_res_57_2,wire_res_57_1,
    wire_res_57_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_29_lo_lo_lo = {wire_res_57_12,wire_res_57_11,wire_res_57_10,wire_res_57_9,wire_res_57_8,
    wire_res_57_7,wire_res_57_6,result_reg_w_29_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_29_lo_lo = {wire_res_57_25,wire_res_57_24,wire_res_57_23,wire_res_57_22,wire_res_57_21,
    wire_res_57_20,wire_res_57_19,result_reg_w_29_lo_lo_hi_lo,result_reg_w_29_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_29_lo = {wire_res_57_52,wire_res_57_51,wire_res_57_50,wire_res_57_49,wire_res_57_48,
    wire_res_57_47,wire_res_57_46,result_reg_w_29_lo_hi_hi_lo,result_reg_w_29_lo_hi_lo,result_reg_w_29_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_29 = {result_reg_w_29_hi,result_reg_w_29_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_58_0 = result_reg_w_29[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_1 = result_reg_w_29[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_2 = result_reg_w_29[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_3 = result_reg_w_29[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_4 = result_reg_w_29[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_5 = result_reg_w_29[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_6 = result_reg_w_29[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_7 = result_reg_w_29[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_8 = result_reg_w_29[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_9 = result_reg_w_29[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_10 = result_reg_w_29[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_11 = result_reg_w_29[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_12 = result_reg_w_29[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_13 = result_reg_w_29[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_14 = result_reg_w_29[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_15 = result_reg_w_29[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_16 = result_reg_w_29[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_17 = result_reg_w_29[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_18 = result_reg_w_29[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_19 = result_reg_w_29[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_20 = result_reg_w_29[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_21 = result_reg_w_29[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_22 = result_reg_w_29[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_23 = result_reg_w_29[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_24 = result_reg_w_29[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_25 = result_reg_w_29[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_26 = result_reg_w_29[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_27 = result_reg_w_29[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_28 = result_reg_w_29[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_29 = result_reg_w_29[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_30 = result_reg_w_29[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_31 = result_reg_w_29[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_32 = result_reg_w_29[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_33 = result_reg_w_29[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_34 = result_reg_w_29[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_35 = result_reg_w_29[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_36 = result_reg_w_29[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_37 = result_reg_w_29[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_38 = result_reg_w_29[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_39 = result_reg_w_29[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_40 = result_reg_w_29[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_41 = result_reg_w_29[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_42 = result_reg_w_29[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_43 = result_reg_w_29[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_44 = result_reg_w_29[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_45 = result_reg_w_29[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_47 = result_reg_w_29[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_48 = result_reg_w_29[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_49 = result_reg_w_29[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_50 = result_reg_w_29[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_51 = result_reg_w_29[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_52 = result_reg_w_29[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_53 = result_reg_w_29[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_54 = result_reg_w_29[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_55 = result_reg_w_29[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_56 = result_reg_w_29[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_57 = result_reg_w_29[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_58 = result_reg_w_29[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_59 = result_reg_w_29[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_60 = result_reg_w_29[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_61 = result_reg_w_29[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_62 = result_reg_w_29[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_63 = result_reg_w_29[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_64 = result_reg_w_29[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_65 = result_reg_w_29[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_66 = result_reg_w_29[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_67 = result_reg_w_29[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_68 = result_reg_w_29[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_69 = result_reg_w_29[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_70 = result_reg_w_29[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_71 = result_reg_w_29[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_72 = result_reg_w_29[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_73 = result_reg_w_29[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_74 = result_reg_w_29[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_75 = result_reg_w_29[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_76 = result_reg_w_29[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_77 = result_reg_w_29[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_78 = result_reg_w_29[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_79 = result_reg_w_29[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_80 = result_reg_w_29[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_81 = result_reg_w_29[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_82 = result_reg_w_29[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_83 = result_reg_w_29[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_84 = result_reg_w_29[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_85 = result_reg_w_29[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_86 = result_reg_w_29[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_87 = result_reg_w_29[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_88 = result_reg_w_29[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_89 = result_reg_w_29[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_90 = result_reg_w_29[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_91 = result_reg_w_29[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_92 = result_reg_w_29[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_93 = result_reg_w_29[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_94 = result_reg_w_29[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_95 = result_reg_w_29[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_96 = result_reg_w_29[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_97 = result_reg_w_29[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_98 = result_reg_w_29[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_99 = result_reg_w_29[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_100 = result_reg_w_29[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_101 = result_reg_w_29[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_102 = result_reg_w_29[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_103 = result_reg_w_29[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_104 = result_reg_w_29[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_58_105 = result_reg_w_29[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_0 = result_reg_r_29[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_1 = result_reg_r_29[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_2 = result_reg_r_29[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_3 = result_reg_r_29[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_4 = result_reg_r_29[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_5 = result_reg_r_29[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_6 = result_reg_r_29[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_7 = result_reg_r_29[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_8 = result_reg_r_29[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_9 = result_reg_r_29[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_10 = result_reg_r_29[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_11 = result_reg_r_29[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_12 = result_reg_r_29[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_13 = result_reg_r_29[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_14 = result_reg_r_29[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_15 = result_reg_r_29[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_16 = result_reg_r_29[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_17 = result_reg_r_29[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_18 = result_reg_r_29[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_19 = result_reg_r_29[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_20 = result_reg_r_29[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_21 = result_reg_r_29[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_22 = result_reg_r_29[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_23 = result_reg_r_29[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_24 = result_reg_r_29[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_25 = result_reg_r_29[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_26 = result_reg_r_29[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_27 = result_reg_r_29[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_28 = result_reg_r_29[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_29 = result_reg_r_29[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_30 = result_reg_r_29[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_31 = result_reg_r_29[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_32 = result_reg_r_29[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_33 = result_reg_r_29[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_34 = result_reg_r_29[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_35 = result_reg_r_29[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_36 = result_reg_r_29[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_37 = result_reg_r_29[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_38 = result_reg_r_29[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_39 = result_reg_r_29[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_40 = result_reg_r_29[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_41 = result_reg_r_29[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_42 = result_reg_r_29[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_43 = result_reg_r_29[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_44 = result_reg_r_29[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_46 = result_reg_r_29[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_47 = result_reg_r_29[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_48 = result_reg_r_29[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_49 = result_reg_r_29[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_50 = result_reg_r_29[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_51 = result_reg_r_29[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_52 = result_reg_r_29[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_53 = result_reg_r_29[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_54 = result_reg_r_29[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_55 = result_reg_r_29[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_56 = result_reg_r_29[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_57 = result_reg_r_29[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_58 = result_reg_r_29[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_59 = result_reg_r_29[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_60 = result_reg_r_29[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_61 = result_reg_r_29[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_62 = result_reg_r_29[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_63 = result_reg_r_29[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_64 = result_reg_r_29[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_65 = result_reg_r_29[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_66 = result_reg_r_29[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_67 = result_reg_r_29[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_68 = result_reg_r_29[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_69 = result_reg_r_29[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_70 = result_reg_r_29[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_71 = result_reg_r_29[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_72 = result_reg_r_29[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_73 = result_reg_r_29[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_74 = result_reg_r_29[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_75 = result_reg_r_29[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_76 = result_reg_r_29[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_77 = result_reg_r_29[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_78 = result_reg_r_29[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_79 = result_reg_r_29[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_80 = result_reg_r_29[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_81 = result_reg_r_29[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_82 = result_reg_r_29[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_83 = result_reg_r_29[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_84 = result_reg_r_29[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_85 = result_reg_r_29[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_86 = result_reg_r_29[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_87 = result_reg_r_29[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_88 = result_reg_r_29[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_89 = result_reg_r_29[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_90 = result_reg_r_29[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_91 = result_reg_r_29[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_92 = result_reg_r_29[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_93 = result_reg_r_29[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_94 = result_reg_r_29[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_95 = result_reg_r_29[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_96 = result_reg_r_29[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_97 = result_reg_r_29[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_98 = result_reg_r_29[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_99 = result_reg_r_29[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_100 = result_reg_r_29[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_101 = result_reg_r_29[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_102 = result_reg_r_29[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_103 = result_reg_r_29[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_104 = result_reg_r_29[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_59_105 = result_reg_r_29[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_30_hi_hi_hi_lo = {wire_res_59_98,wire_res_59_97,wire_res_59_96,wire_res_59_95,wire_res_59_94,
    wire_res_59_93,wire_res_59_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_30_hi_hi_lo_lo = {wire_res_59_84,wire_res_59_83,wire_res_59_82,wire_res_59_81,wire_res_59_80,
    wire_res_59_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_30_hi_hi_lo = {wire_res_59_91,wire_res_59_90,wire_res_59_89,wire_res_59_88,wire_res_59_87,
    wire_res_59_86,wire_res_59_85,result_reg_w_30_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_30_hi_lo_hi_lo = {wire_res_59_71,wire_res_59_70,wire_res_59_69,wire_res_59_68,wire_res_59_67,
    wire_res_59_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_30_hi_lo_lo_lo = {wire_res_59_58,wire_res_59_57,wire_res_59_56,wire_res_59_55,wire_res_59_54,
    wire_res_59_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_30_hi_lo_lo = {wire_res_59_65,wire_res_59_64,wire_res_59_63,wire_res_59_62,wire_res_59_61,
    wire_res_59_60,wire_res_59_59,result_reg_w_30_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_30_hi_lo = {wire_res_59_78,wire_res_59_77,wire_res_59_76,wire_res_59_75,wire_res_59_74,
    wire_res_59_73,wire_res_59_72,result_reg_w_30_hi_lo_hi_lo,result_reg_w_30_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_30_hi = {wire_res_59_105,wire_res_59_104,wire_res_59_103,wire_res_59_102,wire_res_59_101,
    wire_res_59_100,wire_res_59_99,result_reg_w_30_hi_hi_hi_lo,result_reg_w_30_hi_hi_lo,result_reg_w_30_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [150:0] _T_11356 = {b_aux_reg_r_29, 45'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [150:0] _GEN_1301 = {{45'd0}, a_aux_reg_r_29}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_59_45 = _GEN_1301 >= _T_11356; // @[BinaryDesigns2.scala 224:35]
  wire [6:0] result_reg_w_30_lo_hi_hi_lo = {wire_res_59_45,wire_res_59_44,wire_res_59_43,wire_res_59_42,wire_res_59_41,
    wire_res_59_40,wire_res_59_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_30_lo_hi_lo_lo = {wire_res_59_31,wire_res_59_30,wire_res_59_29,wire_res_59_28,wire_res_59_27,
    wire_res_59_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_30_lo_hi_lo = {wire_res_59_38,wire_res_59_37,wire_res_59_36,wire_res_59_35,wire_res_59_34,
    wire_res_59_33,wire_res_59_32,result_reg_w_30_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_30_lo_lo_hi_lo = {wire_res_59_18,wire_res_59_17,wire_res_59_16,wire_res_59_15,wire_res_59_14,
    wire_res_59_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_30_lo_lo_lo_lo = {wire_res_59_5,wire_res_59_4,wire_res_59_3,wire_res_59_2,wire_res_59_1,
    wire_res_59_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_30_lo_lo_lo = {wire_res_59_12,wire_res_59_11,wire_res_59_10,wire_res_59_9,wire_res_59_8,
    wire_res_59_7,wire_res_59_6,result_reg_w_30_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_30_lo_lo = {wire_res_59_25,wire_res_59_24,wire_res_59_23,wire_res_59_22,wire_res_59_21,
    wire_res_59_20,wire_res_59_19,result_reg_w_30_lo_lo_hi_lo,result_reg_w_30_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_30_lo = {wire_res_59_52,wire_res_59_51,wire_res_59_50,wire_res_59_49,wire_res_59_48,
    wire_res_59_47,wire_res_59_46,result_reg_w_30_lo_hi_hi_lo,result_reg_w_30_lo_hi_lo,result_reg_w_30_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_30 = {result_reg_w_30_hi,result_reg_w_30_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_60_0 = result_reg_w_30[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_1 = result_reg_w_30[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_2 = result_reg_w_30[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_3 = result_reg_w_30[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_4 = result_reg_w_30[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_5 = result_reg_w_30[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_6 = result_reg_w_30[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_7 = result_reg_w_30[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_8 = result_reg_w_30[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_9 = result_reg_w_30[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_10 = result_reg_w_30[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_11 = result_reg_w_30[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_12 = result_reg_w_30[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_13 = result_reg_w_30[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_14 = result_reg_w_30[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_15 = result_reg_w_30[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_16 = result_reg_w_30[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_17 = result_reg_w_30[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_18 = result_reg_w_30[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_19 = result_reg_w_30[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_20 = result_reg_w_30[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_21 = result_reg_w_30[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_22 = result_reg_w_30[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_23 = result_reg_w_30[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_24 = result_reg_w_30[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_25 = result_reg_w_30[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_26 = result_reg_w_30[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_27 = result_reg_w_30[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_28 = result_reg_w_30[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_29 = result_reg_w_30[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_30 = result_reg_w_30[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_31 = result_reg_w_30[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_32 = result_reg_w_30[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_33 = result_reg_w_30[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_34 = result_reg_w_30[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_35 = result_reg_w_30[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_36 = result_reg_w_30[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_37 = result_reg_w_30[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_38 = result_reg_w_30[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_39 = result_reg_w_30[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_40 = result_reg_w_30[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_41 = result_reg_w_30[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_42 = result_reg_w_30[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_43 = result_reg_w_30[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_45 = result_reg_w_30[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_46 = result_reg_w_30[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_47 = result_reg_w_30[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_48 = result_reg_w_30[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_49 = result_reg_w_30[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_50 = result_reg_w_30[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_51 = result_reg_w_30[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_52 = result_reg_w_30[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_53 = result_reg_w_30[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_54 = result_reg_w_30[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_55 = result_reg_w_30[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_56 = result_reg_w_30[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_57 = result_reg_w_30[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_58 = result_reg_w_30[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_59 = result_reg_w_30[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_60 = result_reg_w_30[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_61 = result_reg_w_30[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_62 = result_reg_w_30[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_63 = result_reg_w_30[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_64 = result_reg_w_30[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_65 = result_reg_w_30[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_66 = result_reg_w_30[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_67 = result_reg_w_30[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_68 = result_reg_w_30[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_69 = result_reg_w_30[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_70 = result_reg_w_30[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_71 = result_reg_w_30[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_72 = result_reg_w_30[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_73 = result_reg_w_30[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_74 = result_reg_w_30[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_75 = result_reg_w_30[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_76 = result_reg_w_30[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_77 = result_reg_w_30[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_78 = result_reg_w_30[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_79 = result_reg_w_30[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_80 = result_reg_w_30[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_81 = result_reg_w_30[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_82 = result_reg_w_30[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_83 = result_reg_w_30[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_84 = result_reg_w_30[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_85 = result_reg_w_30[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_86 = result_reg_w_30[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_87 = result_reg_w_30[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_88 = result_reg_w_30[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_89 = result_reg_w_30[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_90 = result_reg_w_30[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_91 = result_reg_w_30[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_92 = result_reg_w_30[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_93 = result_reg_w_30[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_94 = result_reg_w_30[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_95 = result_reg_w_30[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_96 = result_reg_w_30[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_97 = result_reg_w_30[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_98 = result_reg_w_30[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_99 = result_reg_w_30[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_100 = result_reg_w_30[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_101 = result_reg_w_30[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_102 = result_reg_w_30[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_103 = result_reg_w_30[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_104 = result_reg_w_30[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_60_105 = result_reg_w_30[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_0 = result_reg_r_30[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_1 = result_reg_r_30[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_2 = result_reg_r_30[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_3 = result_reg_r_30[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_4 = result_reg_r_30[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_5 = result_reg_r_30[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_6 = result_reg_r_30[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_7 = result_reg_r_30[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_8 = result_reg_r_30[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_9 = result_reg_r_30[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_10 = result_reg_r_30[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_11 = result_reg_r_30[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_12 = result_reg_r_30[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_13 = result_reg_r_30[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_14 = result_reg_r_30[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_15 = result_reg_r_30[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_16 = result_reg_r_30[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_17 = result_reg_r_30[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_18 = result_reg_r_30[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_19 = result_reg_r_30[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_20 = result_reg_r_30[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_21 = result_reg_r_30[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_22 = result_reg_r_30[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_23 = result_reg_r_30[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_24 = result_reg_r_30[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_25 = result_reg_r_30[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_26 = result_reg_r_30[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_27 = result_reg_r_30[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_28 = result_reg_r_30[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_29 = result_reg_r_30[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_30 = result_reg_r_30[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_31 = result_reg_r_30[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_32 = result_reg_r_30[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_33 = result_reg_r_30[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_34 = result_reg_r_30[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_35 = result_reg_r_30[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_36 = result_reg_r_30[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_37 = result_reg_r_30[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_38 = result_reg_r_30[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_39 = result_reg_r_30[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_40 = result_reg_r_30[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_41 = result_reg_r_30[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_42 = result_reg_r_30[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_44 = result_reg_r_30[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_45 = result_reg_r_30[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_46 = result_reg_r_30[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_47 = result_reg_r_30[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_48 = result_reg_r_30[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_49 = result_reg_r_30[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_50 = result_reg_r_30[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_51 = result_reg_r_30[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_52 = result_reg_r_30[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_53 = result_reg_r_30[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_54 = result_reg_r_30[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_55 = result_reg_r_30[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_56 = result_reg_r_30[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_57 = result_reg_r_30[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_58 = result_reg_r_30[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_59 = result_reg_r_30[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_60 = result_reg_r_30[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_61 = result_reg_r_30[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_62 = result_reg_r_30[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_63 = result_reg_r_30[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_64 = result_reg_r_30[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_65 = result_reg_r_30[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_66 = result_reg_r_30[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_67 = result_reg_r_30[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_68 = result_reg_r_30[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_69 = result_reg_r_30[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_70 = result_reg_r_30[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_71 = result_reg_r_30[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_72 = result_reg_r_30[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_73 = result_reg_r_30[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_74 = result_reg_r_30[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_75 = result_reg_r_30[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_76 = result_reg_r_30[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_77 = result_reg_r_30[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_78 = result_reg_r_30[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_79 = result_reg_r_30[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_80 = result_reg_r_30[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_81 = result_reg_r_30[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_82 = result_reg_r_30[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_83 = result_reg_r_30[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_84 = result_reg_r_30[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_85 = result_reg_r_30[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_86 = result_reg_r_30[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_87 = result_reg_r_30[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_88 = result_reg_r_30[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_89 = result_reg_r_30[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_90 = result_reg_r_30[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_91 = result_reg_r_30[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_92 = result_reg_r_30[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_93 = result_reg_r_30[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_94 = result_reg_r_30[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_95 = result_reg_r_30[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_96 = result_reg_r_30[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_97 = result_reg_r_30[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_98 = result_reg_r_30[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_99 = result_reg_r_30[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_100 = result_reg_r_30[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_101 = result_reg_r_30[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_102 = result_reg_r_30[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_103 = result_reg_r_30[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_104 = result_reg_r_30[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_61_105 = result_reg_r_30[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_31_hi_hi_hi_lo = {wire_res_61_98,wire_res_61_97,wire_res_61_96,wire_res_61_95,wire_res_61_94,
    wire_res_61_93,wire_res_61_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_31_hi_hi_lo_lo = {wire_res_61_84,wire_res_61_83,wire_res_61_82,wire_res_61_81,wire_res_61_80,
    wire_res_61_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_31_hi_hi_lo = {wire_res_61_91,wire_res_61_90,wire_res_61_89,wire_res_61_88,wire_res_61_87,
    wire_res_61_86,wire_res_61_85,result_reg_w_31_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_31_hi_lo_hi_lo = {wire_res_61_71,wire_res_61_70,wire_res_61_69,wire_res_61_68,wire_res_61_67,
    wire_res_61_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_31_hi_lo_lo_lo = {wire_res_61_58,wire_res_61_57,wire_res_61_56,wire_res_61_55,wire_res_61_54,
    wire_res_61_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_31_hi_lo_lo = {wire_res_61_65,wire_res_61_64,wire_res_61_63,wire_res_61_62,wire_res_61_61,
    wire_res_61_60,wire_res_61_59,result_reg_w_31_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_31_hi_lo = {wire_res_61_78,wire_res_61_77,wire_res_61_76,wire_res_61_75,wire_res_61_74,
    wire_res_61_73,wire_res_61_72,result_reg_w_31_hi_lo_hi_lo,result_reg_w_31_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_31_hi = {wire_res_61_105,wire_res_61_104,wire_res_61_103,wire_res_61_102,wire_res_61_101,
    wire_res_61_100,wire_res_61_99,result_reg_w_31_hi_hi_hi_lo,result_reg_w_31_hi_hi_lo,result_reg_w_31_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [148:0] _T_11360 = {b_aux_reg_r_30, 43'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [148:0] _GEN_1302 = {{43'd0}, a_aux_reg_r_30}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_61_43 = _GEN_1302 >= _T_11360; // @[BinaryDesigns2.scala 224:35]
  wire [6:0] result_reg_w_31_lo_hi_hi_lo = {wire_res_61_45,wire_res_61_44,wire_res_61_43,wire_res_61_42,wire_res_61_41,
    wire_res_61_40,wire_res_61_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_31_lo_hi_lo_lo = {wire_res_61_31,wire_res_61_30,wire_res_61_29,wire_res_61_28,wire_res_61_27,
    wire_res_61_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_31_lo_hi_lo = {wire_res_61_38,wire_res_61_37,wire_res_61_36,wire_res_61_35,wire_res_61_34,
    wire_res_61_33,wire_res_61_32,result_reg_w_31_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_31_lo_lo_hi_lo = {wire_res_61_18,wire_res_61_17,wire_res_61_16,wire_res_61_15,wire_res_61_14,
    wire_res_61_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_31_lo_lo_lo_lo = {wire_res_61_5,wire_res_61_4,wire_res_61_3,wire_res_61_2,wire_res_61_1,
    wire_res_61_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_31_lo_lo_lo = {wire_res_61_12,wire_res_61_11,wire_res_61_10,wire_res_61_9,wire_res_61_8,
    wire_res_61_7,wire_res_61_6,result_reg_w_31_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_31_lo_lo = {wire_res_61_25,wire_res_61_24,wire_res_61_23,wire_res_61_22,wire_res_61_21,
    wire_res_61_20,wire_res_61_19,result_reg_w_31_lo_lo_hi_lo,result_reg_w_31_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_31_lo = {wire_res_61_52,wire_res_61_51,wire_res_61_50,wire_res_61_49,wire_res_61_48,
    wire_res_61_47,wire_res_61_46,result_reg_w_31_lo_hi_hi_lo,result_reg_w_31_lo_hi_lo,result_reg_w_31_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_31 = {result_reg_w_31_hi,result_reg_w_31_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_62_0 = result_reg_w_31[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_1 = result_reg_w_31[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_2 = result_reg_w_31[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_3 = result_reg_w_31[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_4 = result_reg_w_31[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_5 = result_reg_w_31[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_6 = result_reg_w_31[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_7 = result_reg_w_31[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_8 = result_reg_w_31[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_9 = result_reg_w_31[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_10 = result_reg_w_31[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_11 = result_reg_w_31[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_12 = result_reg_w_31[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_13 = result_reg_w_31[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_14 = result_reg_w_31[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_15 = result_reg_w_31[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_16 = result_reg_w_31[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_17 = result_reg_w_31[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_18 = result_reg_w_31[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_19 = result_reg_w_31[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_20 = result_reg_w_31[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_21 = result_reg_w_31[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_22 = result_reg_w_31[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_23 = result_reg_w_31[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_24 = result_reg_w_31[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_25 = result_reg_w_31[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_26 = result_reg_w_31[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_27 = result_reg_w_31[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_28 = result_reg_w_31[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_29 = result_reg_w_31[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_30 = result_reg_w_31[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_31 = result_reg_w_31[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_32 = result_reg_w_31[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_33 = result_reg_w_31[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_34 = result_reg_w_31[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_35 = result_reg_w_31[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_36 = result_reg_w_31[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_37 = result_reg_w_31[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_38 = result_reg_w_31[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_39 = result_reg_w_31[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_40 = result_reg_w_31[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_41 = result_reg_w_31[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_43 = result_reg_w_31[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_44 = result_reg_w_31[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_45 = result_reg_w_31[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_46 = result_reg_w_31[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_47 = result_reg_w_31[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_48 = result_reg_w_31[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_49 = result_reg_w_31[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_50 = result_reg_w_31[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_51 = result_reg_w_31[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_52 = result_reg_w_31[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_53 = result_reg_w_31[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_54 = result_reg_w_31[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_55 = result_reg_w_31[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_56 = result_reg_w_31[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_57 = result_reg_w_31[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_58 = result_reg_w_31[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_59 = result_reg_w_31[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_60 = result_reg_w_31[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_61 = result_reg_w_31[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_62 = result_reg_w_31[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_63 = result_reg_w_31[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_64 = result_reg_w_31[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_65 = result_reg_w_31[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_66 = result_reg_w_31[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_67 = result_reg_w_31[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_68 = result_reg_w_31[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_69 = result_reg_w_31[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_70 = result_reg_w_31[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_71 = result_reg_w_31[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_72 = result_reg_w_31[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_73 = result_reg_w_31[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_74 = result_reg_w_31[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_75 = result_reg_w_31[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_76 = result_reg_w_31[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_77 = result_reg_w_31[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_78 = result_reg_w_31[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_79 = result_reg_w_31[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_80 = result_reg_w_31[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_81 = result_reg_w_31[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_82 = result_reg_w_31[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_83 = result_reg_w_31[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_84 = result_reg_w_31[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_85 = result_reg_w_31[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_86 = result_reg_w_31[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_87 = result_reg_w_31[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_88 = result_reg_w_31[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_89 = result_reg_w_31[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_90 = result_reg_w_31[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_91 = result_reg_w_31[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_92 = result_reg_w_31[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_93 = result_reg_w_31[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_94 = result_reg_w_31[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_95 = result_reg_w_31[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_96 = result_reg_w_31[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_97 = result_reg_w_31[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_98 = result_reg_w_31[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_99 = result_reg_w_31[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_100 = result_reg_w_31[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_101 = result_reg_w_31[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_102 = result_reg_w_31[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_103 = result_reg_w_31[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_104 = result_reg_w_31[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_62_105 = result_reg_w_31[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_0 = result_reg_r_31[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_1 = result_reg_r_31[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_2 = result_reg_r_31[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_3 = result_reg_r_31[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_4 = result_reg_r_31[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_5 = result_reg_r_31[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_6 = result_reg_r_31[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_7 = result_reg_r_31[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_8 = result_reg_r_31[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_9 = result_reg_r_31[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_10 = result_reg_r_31[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_11 = result_reg_r_31[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_12 = result_reg_r_31[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_13 = result_reg_r_31[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_14 = result_reg_r_31[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_15 = result_reg_r_31[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_16 = result_reg_r_31[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_17 = result_reg_r_31[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_18 = result_reg_r_31[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_19 = result_reg_r_31[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_20 = result_reg_r_31[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_21 = result_reg_r_31[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_22 = result_reg_r_31[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_23 = result_reg_r_31[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_24 = result_reg_r_31[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_25 = result_reg_r_31[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_26 = result_reg_r_31[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_27 = result_reg_r_31[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_28 = result_reg_r_31[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_29 = result_reg_r_31[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_30 = result_reg_r_31[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_31 = result_reg_r_31[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_32 = result_reg_r_31[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_33 = result_reg_r_31[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_34 = result_reg_r_31[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_35 = result_reg_r_31[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_36 = result_reg_r_31[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_37 = result_reg_r_31[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_38 = result_reg_r_31[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_39 = result_reg_r_31[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_40 = result_reg_r_31[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_42 = result_reg_r_31[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_43 = result_reg_r_31[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_44 = result_reg_r_31[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_45 = result_reg_r_31[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_46 = result_reg_r_31[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_47 = result_reg_r_31[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_48 = result_reg_r_31[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_49 = result_reg_r_31[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_50 = result_reg_r_31[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_51 = result_reg_r_31[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_52 = result_reg_r_31[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_53 = result_reg_r_31[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_54 = result_reg_r_31[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_55 = result_reg_r_31[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_56 = result_reg_r_31[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_57 = result_reg_r_31[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_58 = result_reg_r_31[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_59 = result_reg_r_31[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_60 = result_reg_r_31[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_61 = result_reg_r_31[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_62 = result_reg_r_31[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_63 = result_reg_r_31[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_64 = result_reg_r_31[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_65 = result_reg_r_31[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_66 = result_reg_r_31[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_67 = result_reg_r_31[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_68 = result_reg_r_31[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_69 = result_reg_r_31[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_70 = result_reg_r_31[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_71 = result_reg_r_31[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_72 = result_reg_r_31[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_73 = result_reg_r_31[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_74 = result_reg_r_31[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_75 = result_reg_r_31[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_76 = result_reg_r_31[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_77 = result_reg_r_31[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_78 = result_reg_r_31[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_79 = result_reg_r_31[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_80 = result_reg_r_31[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_81 = result_reg_r_31[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_82 = result_reg_r_31[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_83 = result_reg_r_31[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_84 = result_reg_r_31[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_85 = result_reg_r_31[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_86 = result_reg_r_31[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_87 = result_reg_r_31[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_88 = result_reg_r_31[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_89 = result_reg_r_31[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_90 = result_reg_r_31[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_91 = result_reg_r_31[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_92 = result_reg_r_31[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_93 = result_reg_r_31[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_94 = result_reg_r_31[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_95 = result_reg_r_31[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_96 = result_reg_r_31[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_97 = result_reg_r_31[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_98 = result_reg_r_31[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_99 = result_reg_r_31[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_100 = result_reg_r_31[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_101 = result_reg_r_31[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_102 = result_reg_r_31[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_103 = result_reg_r_31[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_104 = result_reg_r_31[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_63_105 = result_reg_r_31[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_32_hi_hi_hi_lo = {wire_res_63_98,wire_res_63_97,wire_res_63_96,wire_res_63_95,wire_res_63_94,
    wire_res_63_93,wire_res_63_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_32_hi_hi_lo_lo = {wire_res_63_84,wire_res_63_83,wire_res_63_82,wire_res_63_81,wire_res_63_80,
    wire_res_63_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_32_hi_hi_lo = {wire_res_63_91,wire_res_63_90,wire_res_63_89,wire_res_63_88,wire_res_63_87,
    wire_res_63_86,wire_res_63_85,result_reg_w_32_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_32_hi_lo_hi_lo = {wire_res_63_71,wire_res_63_70,wire_res_63_69,wire_res_63_68,wire_res_63_67,
    wire_res_63_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_32_hi_lo_lo_lo = {wire_res_63_58,wire_res_63_57,wire_res_63_56,wire_res_63_55,wire_res_63_54,
    wire_res_63_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_32_hi_lo_lo = {wire_res_63_65,wire_res_63_64,wire_res_63_63,wire_res_63_62,wire_res_63_61,
    wire_res_63_60,wire_res_63_59,result_reg_w_32_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_32_hi_lo = {wire_res_63_78,wire_res_63_77,wire_res_63_76,wire_res_63_75,wire_res_63_74,
    wire_res_63_73,wire_res_63_72,result_reg_w_32_hi_lo_hi_lo,result_reg_w_32_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_32_hi = {wire_res_63_105,wire_res_63_104,wire_res_63_103,wire_res_63_102,wire_res_63_101,
    wire_res_63_100,wire_res_63_99,result_reg_w_32_hi_hi_hi_lo,result_reg_w_32_hi_hi_lo,result_reg_w_32_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [146:0] _T_11364 = {b_aux_reg_r_31, 41'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [146:0] _GEN_1303 = {{41'd0}, a_aux_reg_r_31}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_63_41 = _GEN_1303 >= _T_11364; // @[BinaryDesigns2.scala 224:35]
  wire [6:0] result_reg_w_32_lo_hi_hi_lo = {wire_res_63_45,wire_res_63_44,wire_res_63_43,wire_res_63_42,wire_res_63_41,
    wire_res_63_40,wire_res_63_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_32_lo_hi_lo_lo = {wire_res_63_31,wire_res_63_30,wire_res_63_29,wire_res_63_28,wire_res_63_27,
    wire_res_63_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_32_lo_hi_lo = {wire_res_63_38,wire_res_63_37,wire_res_63_36,wire_res_63_35,wire_res_63_34,
    wire_res_63_33,wire_res_63_32,result_reg_w_32_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_32_lo_lo_hi_lo = {wire_res_63_18,wire_res_63_17,wire_res_63_16,wire_res_63_15,wire_res_63_14,
    wire_res_63_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_32_lo_lo_lo_lo = {wire_res_63_5,wire_res_63_4,wire_res_63_3,wire_res_63_2,wire_res_63_1,
    wire_res_63_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_32_lo_lo_lo = {wire_res_63_12,wire_res_63_11,wire_res_63_10,wire_res_63_9,wire_res_63_8,
    wire_res_63_7,wire_res_63_6,result_reg_w_32_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_32_lo_lo = {wire_res_63_25,wire_res_63_24,wire_res_63_23,wire_res_63_22,wire_res_63_21,
    wire_res_63_20,wire_res_63_19,result_reg_w_32_lo_lo_hi_lo,result_reg_w_32_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_32_lo = {wire_res_63_52,wire_res_63_51,wire_res_63_50,wire_res_63_49,wire_res_63_48,
    wire_res_63_47,wire_res_63_46,result_reg_w_32_lo_hi_hi_lo,result_reg_w_32_lo_hi_lo,result_reg_w_32_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_32 = {result_reg_w_32_hi,result_reg_w_32_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_64_0 = result_reg_w_32[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_1 = result_reg_w_32[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_2 = result_reg_w_32[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_3 = result_reg_w_32[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_4 = result_reg_w_32[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_5 = result_reg_w_32[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_6 = result_reg_w_32[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_7 = result_reg_w_32[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_8 = result_reg_w_32[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_9 = result_reg_w_32[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_10 = result_reg_w_32[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_11 = result_reg_w_32[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_12 = result_reg_w_32[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_13 = result_reg_w_32[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_14 = result_reg_w_32[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_15 = result_reg_w_32[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_16 = result_reg_w_32[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_17 = result_reg_w_32[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_18 = result_reg_w_32[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_19 = result_reg_w_32[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_20 = result_reg_w_32[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_21 = result_reg_w_32[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_22 = result_reg_w_32[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_23 = result_reg_w_32[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_24 = result_reg_w_32[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_25 = result_reg_w_32[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_26 = result_reg_w_32[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_27 = result_reg_w_32[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_28 = result_reg_w_32[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_29 = result_reg_w_32[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_30 = result_reg_w_32[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_31 = result_reg_w_32[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_32 = result_reg_w_32[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_33 = result_reg_w_32[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_34 = result_reg_w_32[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_35 = result_reg_w_32[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_36 = result_reg_w_32[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_37 = result_reg_w_32[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_38 = result_reg_w_32[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_39 = result_reg_w_32[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_41 = result_reg_w_32[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_42 = result_reg_w_32[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_43 = result_reg_w_32[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_44 = result_reg_w_32[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_45 = result_reg_w_32[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_46 = result_reg_w_32[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_47 = result_reg_w_32[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_48 = result_reg_w_32[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_49 = result_reg_w_32[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_50 = result_reg_w_32[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_51 = result_reg_w_32[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_52 = result_reg_w_32[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_53 = result_reg_w_32[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_54 = result_reg_w_32[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_55 = result_reg_w_32[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_56 = result_reg_w_32[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_57 = result_reg_w_32[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_58 = result_reg_w_32[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_59 = result_reg_w_32[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_60 = result_reg_w_32[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_61 = result_reg_w_32[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_62 = result_reg_w_32[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_63 = result_reg_w_32[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_64 = result_reg_w_32[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_65 = result_reg_w_32[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_66 = result_reg_w_32[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_67 = result_reg_w_32[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_68 = result_reg_w_32[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_69 = result_reg_w_32[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_70 = result_reg_w_32[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_71 = result_reg_w_32[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_72 = result_reg_w_32[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_73 = result_reg_w_32[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_74 = result_reg_w_32[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_75 = result_reg_w_32[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_76 = result_reg_w_32[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_77 = result_reg_w_32[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_78 = result_reg_w_32[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_79 = result_reg_w_32[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_80 = result_reg_w_32[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_81 = result_reg_w_32[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_82 = result_reg_w_32[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_83 = result_reg_w_32[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_84 = result_reg_w_32[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_85 = result_reg_w_32[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_86 = result_reg_w_32[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_87 = result_reg_w_32[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_88 = result_reg_w_32[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_89 = result_reg_w_32[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_90 = result_reg_w_32[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_91 = result_reg_w_32[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_92 = result_reg_w_32[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_93 = result_reg_w_32[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_94 = result_reg_w_32[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_95 = result_reg_w_32[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_96 = result_reg_w_32[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_97 = result_reg_w_32[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_98 = result_reg_w_32[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_99 = result_reg_w_32[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_100 = result_reg_w_32[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_101 = result_reg_w_32[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_102 = result_reg_w_32[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_103 = result_reg_w_32[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_104 = result_reg_w_32[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_64_105 = result_reg_w_32[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_0 = result_reg_r_32[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_1 = result_reg_r_32[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_2 = result_reg_r_32[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_3 = result_reg_r_32[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_4 = result_reg_r_32[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_5 = result_reg_r_32[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_6 = result_reg_r_32[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_7 = result_reg_r_32[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_8 = result_reg_r_32[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_9 = result_reg_r_32[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_10 = result_reg_r_32[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_11 = result_reg_r_32[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_12 = result_reg_r_32[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_13 = result_reg_r_32[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_14 = result_reg_r_32[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_15 = result_reg_r_32[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_16 = result_reg_r_32[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_17 = result_reg_r_32[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_18 = result_reg_r_32[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_19 = result_reg_r_32[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_20 = result_reg_r_32[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_21 = result_reg_r_32[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_22 = result_reg_r_32[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_23 = result_reg_r_32[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_24 = result_reg_r_32[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_25 = result_reg_r_32[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_26 = result_reg_r_32[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_27 = result_reg_r_32[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_28 = result_reg_r_32[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_29 = result_reg_r_32[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_30 = result_reg_r_32[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_31 = result_reg_r_32[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_32 = result_reg_r_32[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_33 = result_reg_r_32[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_34 = result_reg_r_32[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_35 = result_reg_r_32[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_36 = result_reg_r_32[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_37 = result_reg_r_32[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_38 = result_reg_r_32[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_40 = result_reg_r_32[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_41 = result_reg_r_32[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_42 = result_reg_r_32[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_43 = result_reg_r_32[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_44 = result_reg_r_32[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_45 = result_reg_r_32[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_46 = result_reg_r_32[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_47 = result_reg_r_32[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_48 = result_reg_r_32[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_49 = result_reg_r_32[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_50 = result_reg_r_32[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_51 = result_reg_r_32[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_52 = result_reg_r_32[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_53 = result_reg_r_32[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_54 = result_reg_r_32[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_55 = result_reg_r_32[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_56 = result_reg_r_32[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_57 = result_reg_r_32[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_58 = result_reg_r_32[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_59 = result_reg_r_32[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_60 = result_reg_r_32[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_61 = result_reg_r_32[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_62 = result_reg_r_32[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_63 = result_reg_r_32[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_64 = result_reg_r_32[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_65 = result_reg_r_32[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_66 = result_reg_r_32[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_67 = result_reg_r_32[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_68 = result_reg_r_32[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_69 = result_reg_r_32[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_70 = result_reg_r_32[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_71 = result_reg_r_32[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_72 = result_reg_r_32[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_73 = result_reg_r_32[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_74 = result_reg_r_32[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_75 = result_reg_r_32[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_76 = result_reg_r_32[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_77 = result_reg_r_32[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_78 = result_reg_r_32[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_79 = result_reg_r_32[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_80 = result_reg_r_32[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_81 = result_reg_r_32[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_82 = result_reg_r_32[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_83 = result_reg_r_32[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_84 = result_reg_r_32[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_85 = result_reg_r_32[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_86 = result_reg_r_32[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_87 = result_reg_r_32[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_88 = result_reg_r_32[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_89 = result_reg_r_32[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_90 = result_reg_r_32[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_91 = result_reg_r_32[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_92 = result_reg_r_32[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_93 = result_reg_r_32[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_94 = result_reg_r_32[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_95 = result_reg_r_32[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_96 = result_reg_r_32[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_97 = result_reg_r_32[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_98 = result_reg_r_32[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_99 = result_reg_r_32[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_100 = result_reg_r_32[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_101 = result_reg_r_32[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_102 = result_reg_r_32[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_103 = result_reg_r_32[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_104 = result_reg_r_32[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_65_105 = result_reg_r_32[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_33_hi_hi_hi_lo = {wire_res_65_98,wire_res_65_97,wire_res_65_96,wire_res_65_95,wire_res_65_94,
    wire_res_65_93,wire_res_65_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_33_hi_hi_lo_lo = {wire_res_65_84,wire_res_65_83,wire_res_65_82,wire_res_65_81,wire_res_65_80,
    wire_res_65_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_33_hi_hi_lo = {wire_res_65_91,wire_res_65_90,wire_res_65_89,wire_res_65_88,wire_res_65_87,
    wire_res_65_86,wire_res_65_85,result_reg_w_33_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_33_hi_lo_hi_lo = {wire_res_65_71,wire_res_65_70,wire_res_65_69,wire_res_65_68,wire_res_65_67,
    wire_res_65_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_33_hi_lo_lo_lo = {wire_res_65_58,wire_res_65_57,wire_res_65_56,wire_res_65_55,wire_res_65_54,
    wire_res_65_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_33_hi_lo_lo = {wire_res_65_65,wire_res_65_64,wire_res_65_63,wire_res_65_62,wire_res_65_61,
    wire_res_65_60,wire_res_65_59,result_reg_w_33_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_33_hi_lo = {wire_res_65_78,wire_res_65_77,wire_res_65_76,wire_res_65_75,wire_res_65_74,
    wire_res_65_73,wire_res_65_72,result_reg_w_33_hi_lo_hi_lo,result_reg_w_33_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_33_hi = {wire_res_65_105,wire_res_65_104,wire_res_65_103,wire_res_65_102,wire_res_65_101,
    wire_res_65_100,wire_res_65_99,result_reg_w_33_hi_hi_hi_lo,result_reg_w_33_hi_hi_lo,result_reg_w_33_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [144:0] _T_11368 = {b_aux_reg_r_32, 39'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [144:0] _GEN_1304 = {{39'd0}, a_aux_reg_r_32}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_65_39 = _GEN_1304 >= _T_11368; // @[BinaryDesigns2.scala 224:35]
  wire [6:0] result_reg_w_33_lo_hi_hi_lo = {wire_res_65_45,wire_res_65_44,wire_res_65_43,wire_res_65_42,wire_res_65_41,
    wire_res_65_40,wire_res_65_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_33_lo_hi_lo_lo = {wire_res_65_31,wire_res_65_30,wire_res_65_29,wire_res_65_28,wire_res_65_27,
    wire_res_65_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_33_lo_hi_lo = {wire_res_65_38,wire_res_65_37,wire_res_65_36,wire_res_65_35,wire_res_65_34,
    wire_res_65_33,wire_res_65_32,result_reg_w_33_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_33_lo_lo_hi_lo = {wire_res_65_18,wire_res_65_17,wire_res_65_16,wire_res_65_15,wire_res_65_14,
    wire_res_65_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_33_lo_lo_lo_lo = {wire_res_65_5,wire_res_65_4,wire_res_65_3,wire_res_65_2,wire_res_65_1,
    wire_res_65_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_33_lo_lo_lo = {wire_res_65_12,wire_res_65_11,wire_res_65_10,wire_res_65_9,wire_res_65_8,
    wire_res_65_7,wire_res_65_6,result_reg_w_33_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_33_lo_lo = {wire_res_65_25,wire_res_65_24,wire_res_65_23,wire_res_65_22,wire_res_65_21,
    wire_res_65_20,wire_res_65_19,result_reg_w_33_lo_lo_hi_lo,result_reg_w_33_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_33_lo = {wire_res_65_52,wire_res_65_51,wire_res_65_50,wire_res_65_49,wire_res_65_48,
    wire_res_65_47,wire_res_65_46,result_reg_w_33_lo_hi_hi_lo,result_reg_w_33_lo_hi_lo,result_reg_w_33_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_33 = {result_reg_w_33_hi,result_reg_w_33_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_66_0 = result_reg_w_33[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_1 = result_reg_w_33[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_2 = result_reg_w_33[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_3 = result_reg_w_33[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_4 = result_reg_w_33[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_5 = result_reg_w_33[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_6 = result_reg_w_33[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_7 = result_reg_w_33[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_8 = result_reg_w_33[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_9 = result_reg_w_33[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_10 = result_reg_w_33[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_11 = result_reg_w_33[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_12 = result_reg_w_33[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_13 = result_reg_w_33[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_14 = result_reg_w_33[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_15 = result_reg_w_33[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_16 = result_reg_w_33[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_17 = result_reg_w_33[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_18 = result_reg_w_33[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_19 = result_reg_w_33[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_20 = result_reg_w_33[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_21 = result_reg_w_33[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_22 = result_reg_w_33[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_23 = result_reg_w_33[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_24 = result_reg_w_33[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_25 = result_reg_w_33[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_26 = result_reg_w_33[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_27 = result_reg_w_33[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_28 = result_reg_w_33[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_29 = result_reg_w_33[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_30 = result_reg_w_33[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_31 = result_reg_w_33[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_32 = result_reg_w_33[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_33 = result_reg_w_33[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_34 = result_reg_w_33[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_35 = result_reg_w_33[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_36 = result_reg_w_33[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_37 = result_reg_w_33[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_39 = result_reg_w_33[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_40 = result_reg_w_33[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_41 = result_reg_w_33[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_42 = result_reg_w_33[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_43 = result_reg_w_33[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_44 = result_reg_w_33[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_45 = result_reg_w_33[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_46 = result_reg_w_33[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_47 = result_reg_w_33[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_48 = result_reg_w_33[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_49 = result_reg_w_33[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_50 = result_reg_w_33[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_51 = result_reg_w_33[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_52 = result_reg_w_33[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_53 = result_reg_w_33[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_54 = result_reg_w_33[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_55 = result_reg_w_33[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_56 = result_reg_w_33[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_57 = result_reg_w_33[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_58 = result_reg_w_33[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_59 = result_reg_w_33[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_60 = result_reg_w_33[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_61 = result_reg_w_33[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_62 = result_reg_w_33[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_63 = result_reg_w_33[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_64 = result_reg_w_33[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_65 = result_reg_w_33[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_66 = result_reg_w_33[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_67 = result_reg_w_33[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_68 = result_reg_w_33[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_69 = result_reg_w_33[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_70 = result_reg_w_33[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_71 = result_reg_w_33[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_72 = result_reg_w_33[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_73 = result_reg_w_33[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_74 = result_reg_w_33[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_75 = result_reg_w_33[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_76 = result_reg_w_33[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_77 = result_reg_w_33[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_78 = result_reg_w_33[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_79 = result_reg_w_33[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_80 = result_reg_w_33[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_81 = result_reg_w_33[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_82 = result_reg_w_33[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_83 = result_reg_w_33[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_84 = result_reg_w_33[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_85 = result_reg_w_33[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_86 = result_reg_w_33[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_87 = result_reg_w_33[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_88 = result_reg_w_33[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_89 = result_reg_w_33[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_90 = result_reg_w_33[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_91 = result_reg_w_33[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_92 = result_reg_w_33[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_93 = result_reg_w_33[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_94 = result_reg_w_33[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_95 = result_reg_w_33[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_96 = result_reg_w_33[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_97 = result_reg_w_33[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_98 = result_reg_w_33[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_99 = result_reg_w_33[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_100 = result_reg_w_33[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_101 = result_reg_w_33[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_102 = result_reg_w_33[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_103 = result_reg_w_33[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_104 = result_reg_w_33[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_66_105 = result_reg_w_33[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_0 = result_reg_r_33[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_1 = result_reg_r_33[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_2 = result_reg_r_33[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_3 = result_reg_r_33[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_4 = result_reg_r_33[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_5 = result_reg_r_33[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_6 = result_reg_r_33[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_7 = result_reg_r_33[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_8 = result_reg_r_33[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_9 = result_reg_r_33[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_10 = result_reg_r_33[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_11 = result_reg_r_33[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_12 = result_reg_r_33[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_13 = result_reg_r_33[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_14 = result_reg_r_33[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_15 = result_reg_r_33[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_16 = result_reg_r_33[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_17 = result_reg_r_33[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_18 = result_reg_r_33[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_19 = result_reg_r_33[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_20 = result_reg_r_33[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_21 = result_reg_r_33[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_22 = result_reg_r_33[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_23 = result_reg_r_33[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_24 = result_reg_r_33[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_25 = result_reg_r_33[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_26 = result_reg_r_33[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_27 = result_reg_r_33[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_28 = result_reg_r_33[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_29 = result_reg_r_33[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_30 = result_reg_r_33[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_31 = result_reg_r_33[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_32 = result_reg_r_33[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_33 = result_reg_r_33[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_34 = result_reg_r_33[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_35 = result_reg_r_33[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_36 = result_reg_r_33[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_38 = result_reg_r_33[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_39 = result_reg_r_33[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_40 = result_reg_r_33[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_41 = result_reg_r_33[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_42 = result_reg_r_33[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_43 = result_reg_r_33[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_44 = result_reg_r_33[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_45 = result_reg_r_33[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_46 = result_reg_r_33[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_47 = result_reg_r_33[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_48 = result_reg_r_33[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_49 = result_reg_r_33[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_50 = result_reg_r_33[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_51 = result_reg_r_33[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_52 = result_reg_r_33[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_53 = result_reg_r_33[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_54 = result_reg_r_33[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_55 = result_reg_r_33[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_56 = result_reg_r_33[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_57 = result_reg_r_33[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_58 = result_reg_r_33[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_59 = result_reg_r_33[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_60 = result_reg_r_33[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_61 = result_reg_r_33[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_62 = result_reg_r_33[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_63 = result_reg_r_33[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_64 = result_reg_r_33[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_65 = result_reg_r_33[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_66 = result_reg_r_33[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_67 = result_reg_r_33[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_68 = result_reg_r_33[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_69 = result_reg_r_33[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_70 = result_reg_r_33[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_71 = result_reg_r_33[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_72 = result_reg_r_33[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_73 = result_reg_r_33[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_74 = result_reg_r_33[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_75 = result_reg_r_33[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_76 = result_reg_r_33[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_77 = result_reg_r_33[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_78 = result_reg_r_33[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_79 = result_reg_r_33[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_80 = result_reg_r_33[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_81 = result_reg_r_33[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_82 = result_reg_r_33[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_83 = result_reg_r_33[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_84 = result_reg_r_33[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_85 = result_reg_r_33[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_86 = result_reg_r_33[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_87 = result_reg_r_33[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_88 = result_reg_r_33[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_89 = result_reg_r_33[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_90 = result_reg_r_33[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_91 = result_reg_r_33[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_92 = result_reg_r_33[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_93 = result_reg_r_33[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_94 = result_reg_r_33[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_95 = result_reg_r_33[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_96 = result_reg_r_33[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_97 = result_reg_r_33[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_98 = result_reg_r_33[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_99 = result_reg_r_33[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_100 = result_reg_r_33[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_101 = result_reg_r_33[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_102 = result_reg_r_33[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_103 = result_reg_r_33[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_104 = result_reg_r_33[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_67_105 = result_reg_r_33[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_34_hi_hi_hi_lo = {wire_res_67_98,wire_res_67_97,wire_res_67_96,wire_res_67_95,wire_res_67_94,
    wire_res_67_93,wire_res_67_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_34_hi_hi_lo_lo = {wire_res_67_84,wire_res_67_83,wire_res_67_82,wire_res_67_81,wire_res_67_80,
    wire_res_67_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_34_hi_hi_lo = {wire_res_67_91,wire_res_67_90,wire_res_67_89,wire_res_67_88,wire_res_67_87,
    wire_res_67_86,wire_res_67_85,result_reg_w_34_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_34_hi_lo_hi_lo = {wire_res_67_71,wire_res_67_70,wire_res_67_69,wire_res_67_68,wire_res_67_67,
    wire_res_67_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_34_hi_lo_lo_lo = {wire_res_67_58,wire_res_67_57,wire_res_67_56,wire_res_67_55,wire_res_67_54,
    wire_res_67_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_34_hi_lo_lo = {wire_res_67_65,wire_res_67_64,wire_res_67_63,wire_res_67_62,wire_res_67_61,
    wire_res_67_60,wire_res_67_59,result_reg_w_34_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_34_hi_lo = {wire_res_67_78,wire_res_67_77,wire_res_67_76,wire_res_67_75,wire_res_67_74,
    wire_res_67_73,wire_res_67_72,result_reg_w_34_hi_lo_hi_lo,result_reg_w_34_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_34_hi = {wire_res_67_105,wire_res_67_104,wire_res_67_103,wire_res_67_102,wire_res_67_101,
    wire_res_67_100,wire_res_67_99,result_reg_w_34_hi_hi_hi_lo,result_reg_w_34_hi_hi_lo,result_reg_w_34_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_34_lo_hi_hi_lo = {wire_res_67_45,wire_res_67_44,wire_res_67_43,wire_res_67_42,wire_res_67_41,
    wire_res_67_40,wire_res_67_39}; // @[BinaryDesigns2.scala 231:46]
  wire [142:0] _T_11372 = {b_aux_reg_r_33, 37'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [142:0] _GEN_1305 = {{37'd0}, a_aux_reg_r_33}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_67_37 = _GEN_1305 >= _T_11372; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_34_lo_hi_lo_lo = {wire_res_67_31,wire_res_67_30,wire_res_67_29,wire_res_67_28,wire_res_67_27,
    wire_res_67_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_34_lo_hi_lo = {wire_res_67_38,wire_res_67_37,wire_res_67_36,wire_res_67_35,wire_res_67_34,
    wire_res_67_33,wire_res_67_32,result_reg_w_34_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_34_lo_lo_hi_lo = {wire_res_67_18,wire_res_67_17,wire_res_67_16,wire_res_67_15,wire_res_67_14,
    wire_res_67_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_34_lo_lo_lo_lo = {wire_res_67_5,wire_res_67_4,wire_res_67_3,wire_res_67_2,wire_res_67_1,
    wire_res_67_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_34_lo_lo_lo = {wire_res_67_12,wire_res_67_11,wire_res_67_10,wire_res_67_9,wire_res_67_8,
    wire_res_67_7,wire_res_67_6,result_reg_w_34_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_34_lo_lo = {wire_res_67_25,wire_res_67_24,wire_res_67_23,wire_res_67_22,wire_res_67_21,
    wire_res_67_20,wire_res_67_19,result_reg_w_34_lo_lo_hi_lo,result_reg_w_34_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_34_lo = {wire_res_67_52,wire_res_67_51,wire_res_67_50,wire_res_67_49,wire_res_67_48,
    wire_res_67_47,wire_res_67_46,result_reg_w_34_lo_hi_hi_lo,result_reg_w_34_lo_hi_lo,result_reg_w_34_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_34 = {result_reg_w_34_hi,result_reg_w_34_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_68_0 = result_reg_w_34[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_1 = result_reg_w_34[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_2 = result_reg_w_34[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_3 = result_reg_w_34[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_4 = result_reg_w_34[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_5 = result_reg_w_34[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_6 = result_reg_w_34[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_7 = result_reg_w_34[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_8 = result_reg_w_34[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_9 = result_reg_w_34[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_10 = result_reg_w_34[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_11 = result_reg_w_34[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_12 = result_reg_w_34[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_13 = result_reg_w_34[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_14 = result_reg_w_34[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_15 = result_reg_w_34[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_16 = result_reg_w_34[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_17 = result_reg_w_34[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_18 = result_reg_w_34[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_19 = result_reg_w_34[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_20 = result_reg_w_34[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_21 = result_reg_w_34[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_22 = result_reg_w_34[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_23 = result_reg_w_34[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_24 = result_reg_w_34[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_25 = result_reg_w_34[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_26 = result_reg_w_34[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_27 = result_reg_w_34[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_28 = result_reg_w_34[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_29 = result_reg_w_34[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_30 = result_reg_w_34[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_31 = result_reg_w_34[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_32 = result_reg_w_34[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_33 = result_reg_w_34[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_34 = result_reg_w_34[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_35 = result_reg_w_34[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_37 = result_reg_w_34[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_38 = result_reg_w_34[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_39 = result_reg_w_34[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_40 = result_reg_w_34[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_41 = result_reg_w_34[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_42 = result_reg_w_34[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_43 = result_reg_w_34[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_44 = result_reg_w_34[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_45 = result_reg_w_34[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_46 = result_reg_w_34[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_47 = result_reg_w_34[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_48 = result_reg_w_34[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_49 = result_reg_w_34[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_50 = result_reg_w_34[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_51 = result_reg_w_34[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_52 = result_reg_w_34[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_53 = result_reg_w_34[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_54 = result_reg_w_34[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_55 = result_reg_w_34[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_56 = result_reg_w_34[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_57 = result_reg_w_34[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_58 = result_reg_w_34[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_59 = result_reg_w_34[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_60 = result_reg_w_34[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_61 = result_reg_w_34[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_62 = result_reg_w_34[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_63 = result_reg_w_34[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_64 = result_reg_w_34[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_65 = result_reg_w_34[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_66 = result_reg_w_34[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_67 = result_reg_w_34[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_68 = result_reg_w_34[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_69 = result_reg_w_34[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_70 = result_reg_w_34[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_71 = result_reg_w_34[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_72 = result_reg_w_34[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_73 = result_reg_w_34[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_74 = result_reg_w_34[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_75 = result_reg_w_34[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_76 = result_reg_w_34[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_77 = result_reg_w_34[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_78 = result_reg_w_34[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_79 = result_reg_w_34[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_80 = result_reg_w_34[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_81 = result_reg_w_34[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_82 = result_reg_w_34[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_83 = result_reg_w_34[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_84 = result_reg_w_34[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_85 = result_reg_w_34[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_86 = result_reg_w_34[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_87 = result_reg_w_34[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_88 = result_reg_w_34[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_89 = result_reg_w_34[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_90 = result_reg_w_34[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_91 = result_reg_w_34[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_92 = result_reg_w_34[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_93 = result_reg_w_34[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_94 = result_reg_w_34[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_95 = result_reg_w_34[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_96 = result_reg_w_34[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_97 = result_reg_w_34[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_98 = result_reg_w_34[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_99 = result_reg_w_34[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_100 = result_reg_w_34[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_101 = result_reg_w_34[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_102 = result_reg_w_34[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_103 = result_reg_w_34[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_104 = result_reg_w_34[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_68_105 = result_reg_w_34[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_0 = result_reg_r_34[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_1 = result_reg_r_34[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_2 = result_reg_r_34[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_3 = result_reg_r_34[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_4 = result_reg_r_34[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_5 = result_reg_r_34[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_6 = result_reg_r_34[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_7 = result_reg_r_34[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_8 = result_reg_r_34[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_9 = result_reg_r_34[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_10 = result_reg_r_34[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_11 = result_reg_r_34[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_12 = result_reg_r_34[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_13 = result_reg_r_34[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_14 = result_reg_r_34[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_15 = result_reg_r_34[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_16 = result_reg_r_34[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_17 = result_reg_r_34[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_18 = result_reg_r_34[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_19 = result_reg_r_34[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_20 = result_reg_r_34[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_21 = result_reg_r_34[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_22 = result_reg_r_34[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_23 = result_reg_r_34[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_24 = result_reg_r_34[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_25 = result_reg_r_34[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_26 = result_reg_r_34[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_27 = result_reg_r_34[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_28 = result_reg_r_34[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_29 = result_reg_r_34[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_30 = result_reg_r_34[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_31 = result_reg_r_34[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_32 = result_reg_r_34[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_33 = result_reg_r_34[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_34 = result_reg_r_34[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_36 = result_reg_r_34[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_37 = result_reg_r_34[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_38 = result_reg_r_34[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_39 = result_reg_r_34[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_40 = result_reg_r_34[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_41 = result_reg_r_34[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_42 = result_reg_r_34[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_43 = result_reg_r_34[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_44 = result_reg_r_34[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_45 = result_reg_r_34[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_46 = result_reg_r_34[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_47 = result_reg_r_34[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_48 = result_reg_r_34[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_49 = result_reg_r_34[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_50 = result_reg_r_34[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_51 = result_reg_r_34[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_52 = result_reg_r_34[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_53 = result_reg_r_34[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_54 = result_reg_r_34[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_55 = result_reg_r_34[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_56 = result_reg_r_34[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_57 = result_reg_r_34[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_58 = result_reg_r_34[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_59 = result_reg_r_34[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_60 = result_reg_r_34[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_61 = result_reg_r_34[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_62 = result_reg_r_34[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_63 = result_reg_r_34[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_64 = result_reg_r_34[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_65 = result_reg_r_34[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_66 = result_reg_r_34[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_67 = result_reg_r_34[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_68 = result_reg_r_34[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_69 = result_reg_r_34[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_70 = result_reg_r_34[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_71 = result_reg_r_34[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_72 = result_reg_r_34[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_73 = result_reg_r_34[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_74 = result_reg_r_34[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_75 = result_reg_r_34[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_76 = result_reg_r_34[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_77 = result_reg_r_34[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_78 = result_reg_r_34[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_79 = result_reg_r_34[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_80 = result_reg_r_34[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_81 = result_reg_r_34[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_82 = result_reg_r_34[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_83 = result_reg_r_34[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_84 = result_reg_r_34[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_85 = result_reg_r_34[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_86 = result_reg_r_34[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_87 = result_reg_r_34[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_88 = result_reg_r_34[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_89 = result_reg_r_34[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_90 = result_reg_r_34[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_91 = result_reg_r_34[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_92 = result_reg_r_34[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_93 = result_reg_r_34[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_94 = result_reg_r_34[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_95 = result_reg_r_34[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_96 = result_reg_r_34[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_97 = result_reg_r_34[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_98 = result_reg_r_34[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_99 = result_reg_r_34[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_100 = result_reg_r_34[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_101 = result_reg_r_34[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_102 = result_reg_r_34[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_103 = result_reg_r_34[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_104 = result_reg_r_34[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_69_105 = result_reg_r_34[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_35_hi_hi_hi_lo = {wire_res_69_98,wire_res_69_97,wire_res_69_96,wire_res_69_95,wire_res_69_94,
    wire_res_69_93,wire_res_69_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_35_hi_hi_lo_lo = {wire_res_69_84,wire_res_69_83,wire_res_69_82,wire_res_69_81,wire_res_69_80,
    wire_res_69_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_35_hi_hi_lo = {wire_res_69_91,wire_res_69_90,wire_res_69_89,wire_res_69_88,wire_res_69_87,
    wire_res_69_86,wire_res_69_85,result_reg_w_35_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_35_hi_lo_hi_lo = {wire_res_69_71,wire_res_69_70,wire_res_69_69,wire_res_69_68,wire_res_69_67,
    wire_res_69_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_35_hi_lo_lo_lo = {wire_res_69_58,wire_res_69_57,wire_res_69_56,wire_res_69_55,wire_res_69_54,
    wire_res_69_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_35_hi_lo_lo = {wire_res_69_65,wire_res_69_64,wire_res_69_63,wire_res_69_62,wire_res_69_61,
    wire_res_69_60,wire_res_69_59,result_reg_w_35_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_35_hi_lo = {wire_res_69_78,wire_res_69_77,wire_res_69_76,wire_res_69_75,wire_res_69_74,
    wire_res_69_73,wire_res_69_72,result_reg_w_35_hi_lo_hi_lo,result_reg_w_35_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_35_hi = {wire_res_69_105,wire_res_69_104,wire_res_69_103,wire_res_69_102,wire_res_69_101,
    wire_res_69_100,wire_res_69_99,result_reg_w_35_hi_hi_hi_lo,result_reg_w_35_hi_hi_lo,result_reg_w_35_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_35_lo_hi_hi_lo = {wire_res_69_45,wire_res_69_44,wire_res_69_43,wire_res_69_42,wire_res_69_41,
    wire_res_69_40,wire_res_69_39}; // @[BinaryDesigns2.scala 231:46]
  wire [140:0] _T_11376 = {b_aux_reg_r_34, 35'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [140:0] _GEN_1306 = {{35'd0}, a_aux_reg_r_34}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_69_35 = _GEN_1306 >= _T_11376; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_35_lo_hi_lo_lo = {wire_res_69_31,wire_res_69_30,wire_res_69_29,wire_res_69_28,wire_res_69_27,
    wire_res_69_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_35_lo_hi_lo = {wire_res_69_38,wire_res_69_37,wire_res_69_36,wire_res_69_35,wire_res_69_34,
    wire_res_69_33,wire_res_69_32,result_reg_w_35_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_35_lo_lo_hi_lo = {wire_res_69_18,wire_res_69_17,wire_res_69_16,wire_res_69_15,wire_res_69_14,
    wire_res_69_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_35_lo_lo_lo_lo = {wire_res_69_5,wire_res_69_4,wire_res_69_3,wire_res_69_2,wire_res_69_1,
    wire_res_69_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_35_lo_lo_lo = {wire_res_69_12,wire_res_69_11,wire_res_69_10,wire_res_69_9,wire_res_69_8,
    wire_res_69_7,wire_res_69_6,result_reg_w_35_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_35_lo_lo = {wire_res_69_25,wire_res_69_24,wire_res_69_23,wire_res_69_22,wire_res_69_21,
    wire_res_69_20,wire_res_69_19,result_reg_w_35_lo_lo_hi_lo,result_reg_w_35_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_35_lo = {wire_res_69_52,wire_res_69_51,wire_res_69_50,wire_res_69_49,wire_res_69_48,
    wire_res_69_47,wire_res_69_46,result_reg_w_35_lo_hi_hi_lo,result_reg_w_35_lo_hi_lo,result_reg_w_35_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_35 = {result_reg_w_35_hi,result_reg_w_35_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_70_0 = result_reg_w_35[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_1 = result_reg_w_35[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_2 = result_reg_w_35[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_3 = result_reg_w_35[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_4 = result_reg_w_35[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_5 = result_reg_w_35[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_6 = result_reg_w_35[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_7 = result_reg_w_35[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_8 = result_reg_w_35[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_9 = result_reg_w_35[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_10 = result_reg_w_35[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_11 = result_reg_w_35[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_12 = result_reg_w_35[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_13 = result_reg_w_35[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_14 = result_reg_w_35[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_15 = result_reg_w_35[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_16 = result_reg_w_35[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_17 = result_reg_w_35[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_18 = result_reg_w_35[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_19 = result_reg_w_35[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_20 = result_reg_w_35[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_21 = result_reg_w_35[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_22 = result_reg_w_35[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_23 = result_reg_w_35[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_24 = result_reg_w_35[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_25 = result_reg_w_35[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_26 = result_reg_w_35[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_27 = result_reg_w_35[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_28 = result_reg_w_35[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_29 = result_reg_w_35[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_30 = result_reg_w_35[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_31 = result_reg_w_35[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_32 = result_reg_w_35[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_33 = result_reg_w_35[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_35 = result_reg_w_35[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_36 = result_reg_w_35[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_37 = result_reg_w_35[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_38 = result_reg_w_35[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_39 = result_reg_w_35[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_40 = result_reg_w_35[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_41 = result_reg_w_35[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_42 = result_reg_w_35[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_43 = result_reg_w_35[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_44 = result_reg_w_35[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_45 = result_reg_w_35[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_46 = result_reg_w_35[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_47 = result_reg_w_35[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_48 = result_reg_w_35[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_49 = result_reg_w_35[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_50 = result_reg_w_35[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_51 = result_reg_w_35[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_52 = result_reg_w_35[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_53 = result_reg_w_35[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_54 = result_reg_w_35[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_55 = result_reg_w_35[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_56 = result_reg_w_35[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_57 = result_reg_w_35[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_58 = result_reg_w_35[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_59 = result_reg_w_35[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_60 = result_reg_w_35[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_61 = result_reg_w_35[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_62 = result_reg_w_35[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_63 = result_reg_w_35[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_64 = result_reg_w_35[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_65 = result_reg_w_35[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_66 = result_reg_w_35[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_67 = result_reg_w_35[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_68 = result_reg_w_35[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_69 = result_reg_w_35[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_70 = result_reg_w_35[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_71 = result_reg_w_35[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_72 = result_reg_w_35[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_73 = result_reg_w_35[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_74 = result_reg_w_35[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_75 = result_reg_w_35[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_76 = result_reg_w_35[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_77 = result_reg_w_35[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_78 = result_reg_w_35[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_79 = result_reg_w_35[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_80 = result_reg_w_35[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_81 = result_reg_w_35[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_82 = result_reg_w_35[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_83 = result_reg_w_35[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_84 = result_reg_w_35[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_85 = result_reg_w_35[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_86 = result_reg_w_35[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_87 = result_reg_w_35[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_88 = result_reg_w_35[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_89 = result_reg_w_35[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_90 = result_reg_w_35[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_91 = result_reg_w_35[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_92 = result_reg_w_35[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_93 = result_reg_w_35[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_94 = result_reg_w_35[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_95 = result_reg_w_35[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_96 = result_reg_w_35[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_97 = result_reg_w_35[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_98 = result_reg_w_35[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_99 = result_reg_w_35[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_100 = result_reg_w_35[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_101 = result_reg_w_35[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_102 = result_reg_w_35[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_103 = result_reg_w_35[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_104 = result_reg_w_35[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_70_105 = result_reg_w_35[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_0 = result_reg_r_35[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_1 = result_reg_r_35[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_2 = result_reg_r_35[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_3 = result_reg_r_35[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_4 = result_reg_r_35[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_5 = result_reg_r_35[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_6 = result_reg_r_35[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_7 = result_reg_r_35[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_8 = result_reg_r_35[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_9 = result_reg_r_35[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_10 = result_reg_r_35[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_11 = result_reg_r_35[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_12 = result_reg_r_35[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_13 = result_reg_r_35[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_14 = result_reg_r_35[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_15 = result_reg_r_35[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_16 = result_reg_r_35[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_17 = result_reg_r_35[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_18 = result_reg_r_35[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_19 = result_reg_r_35[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_20 = result_reg_r_35[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_21 = result_reg_r_35[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_22 = result_reg_r_35[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_23 = result_reg_r_35[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_24 = result_reg_r_35[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_25 = result_reg_r_35[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_26 = result_reg_r_35[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_27 = result_reg_r_35[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_28 = result_reg_r_35[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_29 = result_reg_r_35[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_30 = result_reg_r_35[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_31 = result_reg_r_35[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_32 = result_reg_r_35[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_34 = result_reg_r_35[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_35 = result_reg_r_35[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_36 = result_reg_r_35[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_37 = result_reg_r_35[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_38 = result_reg_r_35[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_39 = result_reg_r_35[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_40 = result_reg_r_35[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_41 = result_reg_r_35[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_42 = result_reg_r_35[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_43 = result_reg_r_35[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_44 = result_reg_r_35[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_45 = result_reg_r_35[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_46 = result_reg_r_35[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_47 = result_reg_r_35[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_48 = result_reg_r_35[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_49 = result_reg_r_35[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_50 = result_reg_r_35[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_51 = result_reg_r_35[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_52 = result_reg_r_35[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_53 = result_reg_r_35[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_54 = result_reg_r_35[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_55 = result_reg_r_35[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_56 = result_reg_r_35[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_57 = result_reg_r_35[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_58 = result_reg_r_35[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_59 = result_reg_r_35[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_60 = result_reg_r_35[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_61 = result_reg_r_35[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_62 = result_reg_r_35[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_63 = result_reg_r_35[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_64 = result_reg_r_35[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_65 = result_reg_r_35[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_66 = result_reg_r_35[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_67 = result_reg_r_35[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_68 = result_reg_r_35[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_69 = result_reg_r_35[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_70 = result_reg_r_35[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_71 = result_reg_r_35[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_72 = result_reg_r_35[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_73 = result_reg_r_35[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_74 = result_reg_r_35[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_75 = result_reg_r_35[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_76 = result_reg_r_35[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_77 = result_reg_r_35[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_78 = result_reg_r_35[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_79 = result_reg_r_35[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_80 = result_reg_r_35[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_81 = result_reg_r_35[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_82 = result_reg_r_35[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_83 = result_reg_r_35[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_84 = result_reg_r_35[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_85 = result_reg_r_35[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_86 = result_reg_r_35[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_87 = result_reg_r_35[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_88 = result_reg_r_35[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_89 = result_reg_r_35[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_90 = result_reg_r_35[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_91 = result_reg_r_35[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_92 = result_reg_r_35[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_93 = result_reg_r_35[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_94 = result_reg_r_35[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_95 = result_reg_r_35[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_96 = result_reg_r_35[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_97 = result_reg_r_35[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_98 = result_reg_r_35[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_99 = result_reg_r_35[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_100 = result_reg_r_35[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_101 = result_reg_r_35[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_102 = result_reg_r_35[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_103 = result_reg_r_35[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_104 = result_reg_r_35[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_71_105 = result_reg_r_35[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_36_hi_hi_hi_lo = {wire_res_71_98,wire_res_71_97,wire_res_71_96,wire_res_71_95,wire_res_71_94,
    wire_res_71_93,wire_res_71_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_36_hi_hi_lo_lo = {wire_res_71_84,wire_res_71_83,wire_res_71_82,wire_res_71_81,wire_res_71_80,
    wire_res_71_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_36_hi_hi_lo = {wire_res_71_91,wire_res_71_90,wire_res_71_89,wire_res_71_88,wire_res_71_87,
    wire_res_71_86,wire_res_71_85,result_reg_w_36_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_36_hi_lo_hi_lo = {wire_res_71_71,wire_res_71_70,wire_res_71_69,wire_res_71_68,wire_res_71_67,
    wire_res_71_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_36_hi_lo_lo_lo = {wire_res_71_58,wire_res_71_57,wire_res_71_56,wire_res_71_55,wire_res_71_54,
    wire_res_71_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_36_hi_lo_lo = {wire_res_71_65,wire_res_71_64,wire_res_71_63,wire_res_71_62,wire_res_71_61,
    wire_res_71_60,wire_res_71_59,result_reg_w_36_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_36_hi_lo = {wire_res_71_78,wire_res_71_77,wire_res_71_76,wire_res_71_75,wire_res_71_74,
    wire_res_71_73,wire_res_71_72,result_reg_w_36_hi_lo_hi_lo,result_reg_w_36_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_36_hi = {wire_res_71_105,wire_res_71_104,wire_res_71_103,wire_res_71_102,wire_res_71_101,
    wire_res_71_100,wire_res_71_99,result_reg_w_36_hi_hi_hi_lo,result_reg_w_36_hi_hi_lo,result_reg_w_36_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_36_lo_hi_hi_lo = {wire_res_71_45,wire_res_71_44,wire_res_71_43,wire_res_71_42,wire_res_71_41,
    wire_res_71_40,wire_res_71_39}; // @[BinaryDesigns2.scala 231:46]
  wire [138:0] _T_11380 = {b_aux_reg_r_35, 33'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [138:0] _GEN_1307 = {{33'd0}, a_aux_reg_r_35}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_71_33 = _GEN_1307 >= _T_11380; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_36_lo_hi_lo_lo = {wire_res_71_31,wire_res_71_30,wire_res_71_29,wire_res_71_28,wire_res_71_27,
    wire_res_71_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_36_lo_hi_lo = {wire_res_71_38,wire_res_71_37,wire_res_71_36,wire_res_71_35,wire_res_71_34,
    wire_res_71_33,wire_res_71_32,result_reg_w_36_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_36_lo_lo_hi_lo = {wire_res_71_18,wire_res_71_17,wire_res_71_16,wire_res_71_15,wire_res_71_14,
    wire_res_71_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_36_lo_lo_lo_lo = {wire_res_71_5,wire_res_71_4,wire_res_71_3,wire_res_71_2,wire_res_71_1,
    wire_res_71_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_36_lo_lo_lo = {wire_res_71_12,wire_res_71_11,wire_res_71_10,wire_res_71_9,wire_res_71_8,
    wire_res_71_7,wire_res_71_6,result_reg_w_36_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_36_lo_lo = {wire_res_71_25,wire_res_71_24,wire_res_71_23,wire_res_71_22,wire_res_71_21,
    wire_res_71_20,wire_res_71_19,result_reg_w_36_lo_lo_hi_lo,result_reg_w_36_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_36_lo = {wire_res_71_52,wire_res_71_51,wire_res_71_50,wire_res_71_49,wire_res_71_48,
    wire_res_71_47,wire_res_71_46,result_reg_w_36_lo_hi_hi_lo,result_reg_w_36_lo_hi_lo,result_reg_w_36_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_36 = {result_reg_w_36_hi,result_reg_w_36_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_72_0 = result_reg_w_36[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_1 = result_reg_w_36[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_2 = result_reg_w_36[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_3 = result_reg_w_36[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_4 = result_reg_w_36[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_5 = result_reg_w_36[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_6 = result_reg_w_36[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_7 = result_reg_w_36[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_8 = result_reg_w_36[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_9 = result_reg_w_36[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_10 = result_reg_w_36[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_11 = result_reg_w_36[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_12 = result_reg_w_36[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_13 = result_reg_w_36[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_14 = result_reg_w_36[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_15 = result_reg_w_36[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_16 = result_reg_w_36[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_17 = result_reg_w_36[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_18 = result_reg_w_36[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_19 = result_reg_w_36[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_20 = result_reg_w_36[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_21 = result_reg_w_36[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_22 = result_reg_w_36[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_23 = result_reg_w_36[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_24 = result_reg_w_36[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_25 = result_reg_w_36[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_26 = result_reg_w_36[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_27 = result_reg_w_36[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_28 = result_reg_w_36[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_29 = result_reg_w_36[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_30 = result_reg_w_36[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_31 = result_reg_w_36[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_33 = result_reg_w_36[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_34 = result_reg_w_36[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_35 = result_reg_w_36[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_36 = result_reg_w_36[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_37 = result_reg_w_36[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_38 = result_reg_w_36[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_39 = result_reg_w_36[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_40 = result_reg_w_36[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_41 = result_reg_w_36[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_42 = result_reg_w_36[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_43 = result_reg_w_36[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_44 = result_reg_w_36[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_45 = result_reg_w_36[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_46 = result_reg_w_36[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_47 = result_reg_w_36[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_48 = result_reg_w_36[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_49 = result_reg_w_36[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_50 = result_reg_w_36[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_51 = result_reg_w_36[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_52 = result_reg_w_36[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_53 = result_reg_w_36[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_54 = result_reg_w_36[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_55 = result_reg_w_36[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_56 = result_reg_w_36[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_57 = result_reg_w_36[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_58 = result_reg_w_36[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_59 = result_reg_w_36[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_60 = result_reg_w_36[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_61 = result_reg_w_36[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_62 = result_reg_w_36[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_63 = result_reg_w_36[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_64 = result_reg_w_36[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_65 = result_reg_w_36[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_66 = result_reg_w_36[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_67 = result_reg_w_36[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_68 = result_reg_w_36[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_69 = result_reg_w_36[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_70 = result_reg_w_36[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_71 = result_reg_w_36[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_72 = result_reg_w_36[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_73 = result_reg_w_36[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_74 = result_reg_w_36[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_75 = result_reg_w_36[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_76 = result_reg_w_36[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_77 = result_reg_w_36[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_78 = result_reg_w_36[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_79 = result_reg_w_36[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_80 = result_reg_w_36[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_81 = result_reg_w_36[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_82 = result_reg_w_36[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_83 = result_reg_w_36[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_84 = result_reg_w_36[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_85 = result_reg_w_36[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_86 = result_reg_w_36[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_87 = result_reg_w_36[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_88 = result_reg_w_36[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_89 = result_reg_w_36[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_90 = result_reg_w_36[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_91 = result_reg_w_36[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_92 = result_reg_w_36[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_93 = result_reg_w_36[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_94 = result_reg_w_36[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_95 = result_reg_w_36[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_96 = result_reg_w_36[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_97 = result_reg_w_36[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_98 = result_reg_w_36[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_99 = result_reg_w_36[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_100 = result_reg_w_36[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_101 = result_reg_w_36[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_102 = result_reg_w_36[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_103 = result_reg_w_36[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_104 = result_reg_w_36[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_72_105 = result_reg_w_36[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_0 = result_reg_r_36[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_1 = result_reg_r_36[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_2 = result_reg_r_36[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_3 = result_reg_r_36[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_4 = result_reg_r_36[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_5 = result_reg_r_36[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_6 = result_reg_r_36[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_7 = result_reg_r_36[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_8 = result_reg_r_36[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_9 = result_reg_r_36[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_10 = result_reg_r_36[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_11 = result_reg_r_36[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_12 = result_reg_r_36[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_13 = result_reg_r_36[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_14 = result_reg_r_36[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_15 = result_reg_r_36[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_16 = result_reg_r_36[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_17 = result_reg_r_36[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_18 = result_reg_r_36[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_19 = result_reg_r_36[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_20 = result_reg_r_36[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_21 = result_reg_r_36[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_22 = result_reg_r_36[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_23 = result_reg_r_36[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_24 = result_reg_r_36[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_25 = result_reg_r_36[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_26 = result_reg_r_36[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_27 = result_reg_r_36[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_28 = result_reg_r_36[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_29 = result_reg_r_36[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_30 = result_reg_r_36[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_32 = result_reg_r_36[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_33 = result_reg_r_36[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_34 = result_reg_r_36[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_35 = result_reg_r_36[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_36 = result_reg_r_36[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_37 = result_reg_r_36[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_38 = result_reg_r_36[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_39 = result_reg_r_36[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_40 = result_reg_r_36[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_41 = result_reg_r_36[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_42 = result_reg_r_36[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_43 = result_reg_r_36[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_44 = result_reg_r_36[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_45 = result_reg_r_36[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_46 = result_reg_r_36[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_47 = result_reg_r_36[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_48 = result_reg_r_36[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_49 = result_reg_r_36[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_50 = result_reg_r_36[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_51 = result_reg_r_36[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_52 = result_reg_r_36[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_53 = result_reg_r_36[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_54 = result_reg_r_36[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_55 = result_reg_r_36[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_56 = result_reg_r_36[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_57 = result_reg_r_36[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_58 = result_reg_r_36[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_59 = result_reg_r_36[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_60 = result_reg_r_36[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_61 = result_reg_r_36[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_62 = result_reg_r_36[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_63 = result_reg_r_36[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_64 = result_reg_r_36[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_65 = result_reg_r_36[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_66 = result_reg_r_36[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_67 = result_reg_r_36[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_68 = result_reg_r_36[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_69 = result_reg_r_36[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_70 = result_reg_r_36[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_71 = result_reg_r_36[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_72 = result_reg_r_36[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_73 = result_reg_r_36[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_74 = result_reg_r_36[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_75 = result_reg_r_36[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_76 = result_reg_r_36[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_77 = result_reg_r_36[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_78 = result_reg_r_36[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_79 = result_reg_r_36[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_80 = result_reg_r_36[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_81 = result_reg_r_36[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_82 = result_reg_r_36[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_83 = result_reg_r_36[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_84 = result_reg_r_36[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_85 = result_reg_r_36[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_86 = result_reg_r_36[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_87 = result_reg_r_36[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_88 = result_reg_r_36[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_89 = result_reg_r_36[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_90 = result_reg_r_36[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_91 = result_reg_r_36[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_92 = result_reg_r_36[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_93 = result_reg_r_36[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_94 = result_reg_r_36[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_95 = result_reg_r_36[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_96 = result_reg_r_36[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_97 = result_reg_r_36[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_98 = result_reg_r_36[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_99 = result_reg_r_36[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_100 = result_reg_r_36[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_101 = result_reg_r_36[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_102 = result_reg_r_36[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_103 = result_reg_r_36[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_104 = result_reg_r_36[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_73_105 = result_reg_r_36[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_37_hi_hi_hi_lo = {wire_res_73_98,wire_res_73_97,wire_res_73_96,wire_res_73_95,wire_res_73_94,
    wire_res_73_93,wire_res_73_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_37_hi_hi_lo_lo = {wire_res_73_84,wire_res_73_83,wire_res_73_82,wire_res_73_81,wire_res_73_80,
    wire_res_73_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_37_hi_hi_lo = {wire_res_73_91,wire_res_73_90,wire_res_73_89,wire_res_73_88,wire_res_73_87,
    wire_res_73_86,wire_res_73_85,result_reg_w_37_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_37_hi_lo_hi_lo = {wire_res_73_71,wire_res_73_70,wire_res_73_69,wire_res_73_68,wire_res_73_67,
    wire_res_73_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_37_hi_lo_lo_lo = {wire_res_73_58,wire_res_73_57,wire_res_73_56,wire_res_73_55,wire_res_73_54,
    wire_res_73_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_37_hi_lo_lo = {wire_res_73_65,wire_res_73_64,wire_res_73_63,wire_res_73_62,wire_res_73_61,
    wire_res_73_60,wire_res_73_59,result_reg_w_37_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_37_hi_lo = {wire_res_73_78,wire_res_73_77,wire_res_73_76,wire_res_73_75,wire_res_73_74,
    wire_res_73_73,wire_res_73_72,result_reg_w_37_hi_lo_hi_lo,result_reg_w_37_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_37_hi = {wire_res_73_105,wire_res_73_104,wire_res_73_103,wire_res_73_102,wire_res_73_101,
    wire_res_73_100,wire_res_73_99,result_reg_w_37_hi_hi_hi_lo,result_reg_w_37_hi_hi_lo,result_reg_w_37_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_37_lo_hi_hi_lo = {wire_res_73_45,wire_res_73_44,wire_res_73_43,wire_res_73_42,wire_res_73_41,
    wire_res_73_40,wire_res_73_39}; // @[BinaryDesigns2.scala 231:46]
  wire [136:0] _T_11384 = {b_aux_reg_r_36, 31'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [136:0] _GEN_1308 = {{31'd0}, a_aux_reg_r_36}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_73_31 = _GEN_1308 >= _T_11384; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_37_lo_hi_lo_lo = {wire_res_73_31,wire_res_73_30,wire_res_73_29,wire_res_73_28,wire_res_73_27,
    wire_res_73_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_37_lo_hi_lo = {wire_res_73_38,wire_res_73_37,wire_res_73_36,wire_res_73_35,wire_res_73_34,
    wire_res_73_33,wire_res_73_32,result_reg_w_37_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_37_lo_lo_hi_lo = {wire_res_73_18,wire_res_73_17,wire_res_73_16,wire_res_73_15,wire_res_73_14,
    wire_res_73_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_37_lo_lo_lo_lo = {wire_res_73_5,wire_res_73_4,wire_res_73_3,wire_res_73_2,wire_res_73_1,
    wire_res_73_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_37_lo_lo_lo = {wire_res_73_12,wire_res_73_11,wire_res_73_10,wire_res_73_9,wire_res_73_8,
    wire_res_73_7,wire_res_73_6,result_reg_w_37_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_37_lo_lo = {wire_res_73_25,wire_res_73_24,wire_res_73_23,wire_res_73_22,wire_res_73_21,
    wire_res_73_20,wire_res_73_19,result_reg_w_37_lo_lo_hi_lo,result_reg_w_37_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_37_lo = {wire_res_73_52,wire_res_73_51,wire_res_73_50,wire_res_73_49,wire_res_73_48,
    wire_res_73_47,wire_res_73_46,result_reg_w_37_lo_hi_hi_lo,result_reg_w_37_lo_hi_lo,result_reg_w_37_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_37 = {result_reg_w_37_hi,result_reg_w_37_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_74_0 = result_reg_w_37[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_1 = result_reg_w_37[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_2 = result_reg_w_37[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_3 = result_reg_w_37[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_4 = result_reg_w_37[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_5 = result_reg_w_37[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_6 = result_reg_w_37[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_7 = result_reg_w_37[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_8 = result_reg_w_37[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_9 = result_reg_w_37[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_10 = result_reg_w_37[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_11 = result_reg_w_37[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_12 = result_reg_w_37[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_13 = result_reg_w_37[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_14 = result_reg_w_37[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_15 = result_reg_w_37[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_16 = result_reg_w_37[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_17 = result_reg_w_37[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_18 = result_reg_w_37[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_19 = result_reg_w_37[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_20 = result_reg_w_37[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_21 = result_reg_w_37[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_22 = result_reg_w_37[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_23 = result_reg_w_37[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_24 = result_reg_w_37[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_25 = result_reg_w_37[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_26 = result_reg_w_37[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_27 = result_reg_w_37[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_28 = result_reg_w_37[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_29 = result_reg_w_37[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_31 = result_reg_w_37[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_32 = result_reg_w_37[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_33 = result_reg_w_37[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_34 = result_reg_w_37[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_35 = result_reg_w_37[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_36 = result_reg_w_37[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_37 = result_reg_w_37[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_38 = result_reg_w_37[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_39 = result_reg_w_37[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_40 = result_reg_w_37[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_41 = result_reg_w_37[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_42 = result_reg_w_37[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_43 = result_reg_w_37[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_44 = result_reg_w_37[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_45 = result_reg_w_37[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_46 = result_reg_w_37[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_47 = result_reg_w_37[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_48 = result_reg_w_37[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_49 = result_reg_w_37[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_50 = result_reg_w_37[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_51 = result_reg_w_37[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_52 = result_reg_w_37[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_53 = result_reg_w_37[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_54 = result_reg_w_37[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_55 = result_reg_w_37[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_56 = result_reg_w_37[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_57 = result_reg_w_37[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_58 = result_reg_w_37[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_59 = result_reg_w_37[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_60 = result_reg_w_37[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_61 = result_reg_w_37[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_62 = result_reg_w_37[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_63 = result_reg_w_37[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_64 = result_reg_w_37[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_65 = result_reg_w_37[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_66 = result_reg_w_37[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_67 = result_reg_w_37[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_68 = result_reg_w_37[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_69 = result_reg_w_37[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_70 = result_reg_w_37[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_71 = result_reg_w_37[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_72 = result_reg_w_37[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_73 = result_reg_w_37[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_74 = result_reg_w_37[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_75 = result_reg_w_37[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_76 = result_reg_w_37[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_77 = result_reg_w_37[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_78 = result_reg_w_37[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_79 = result_reg_w_37[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_80 = result_reg_w_37[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_81 = result_reg_w_37[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_82 = result_reg_w_37[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_83 = result_reg_w_37[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_84 = result_reg_w_37[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_85 = result_reg_w_37[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_86 = result_reg_w_37[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_87 = result_reg_w_37[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_88 = result_reg_w_37[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_89 = result_reg_w_37[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_90 = result_reg_w_37[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_91 = result_reg_w_37[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_92 = result_reg_w_37[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_93 = result_reg_w_37[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_94 = result_reg_w_37[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_95 = result_reg_w_37[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_96 = result_reg_w_37[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_97 = result_reg_w_37[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_98 = result_reg_w_37[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_99 = result_reg_w_37[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_100 = result_reg_w_37[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_101 = result_reg_w_37[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_102 = result_reg_w_37[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_103 = result_reg_w_37[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_104 = result_reg_w_37[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_74_105 = result_reg_w_37[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_0 = result_reg_r_37[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_1 = result_reg_r_37[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_2 = result_reg_r_37[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_3 = result_reg_r_37[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_4 = result_reg_r_37[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_5 = result_reg_r_37[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_6 = result_reg_r_37[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_7 = result_reg_r_37[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_8 = result_reg_r_37[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_9 = result_reg_r_37[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_10 = result_reg_r_37[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_11 = result_reg_r_37[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_12 = result_reg_r_37[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_13 = result_reg_r_37[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_14 = result_reg_r_37[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_15 = result_reg_r_37[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_16 = result_reg_r_37[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_17 = result_reg_r_37[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_18 = result_reg_r_37[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_19 = result_reg_r_37[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_20 = result_reg_r_37[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_21 = result_reg_r_37[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_22 = result_reg_r_37[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_23 = result_reg_r_37[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_24 = result_reg_r_37[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_25 = result_reg_r_37[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_26 = result_reg_r_37[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_27 = result_reg_r_37[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_28 = result_reg_r_37[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_30 = result_reg_r_37[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_31 = result_reg_r_37[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_32 = result_reg_r_37[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_33 = result_reg_r_37[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_34 = result_reg_r_37[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_35 = result_reg_r_37[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_36 = result_reg_r_37[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_37 = result_reg_r_37[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_38 = result_reg_r_37[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_39 = result_reg_r_37[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_40 = result_reg_r_37[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_41 = result_reg_r_37[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_42 = result_reg_r_37[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_43 = result_reg_r_37[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_44 = result_reg_r_37[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_45 = result_reg_r_37[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_46 = result_reg_r_37[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_47 = result_reg_r_37[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_48 = result_reg_r_37[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_49 = result_reg_r_37[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_50 = result_reg_r_37[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_51 = result_reg_r_37[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_52 = result_reg_r_37[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_53 = result_reg_r_37[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_54 = result_reg_r_37[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_55 = result_reg_r_37[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_56 = result_reg_r_37[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_57 = result_reg_r_37[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_58 = result_reg_r_37[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_59 = result_reg_r_37[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_60 = result_reg_r_37[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_61 = result_reg_r_37[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_62 = result_reg_r_37[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_63 = result_reg_r_37[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_64 = result_reg_r_37[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_65 = result_reg_r_37[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_66 = result_reg_r_37[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_67 = result_reg_r_37[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_68 = result_reg_r_37[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_69 = result_reg_r_37[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_70 = result_reg_r_37[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_71 = result_reg_r_37[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_72 = result_reg_r_37[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_73 = result_reg_r_37[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_74 = result_reg_r_37[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_75 = result_reg_r_37[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_76 = result_reg_r_37[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_77 = result_reg_r_37[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_78 = result_reg_r_37[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_79 = result_reg_r_37[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_80 = result_reg_r_37[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_81 = result_reg_r_37[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_82 = result_reg_r_37[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_83 = result_reg_r_37[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_84 = result_reg_r_37[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_85 = result_reg_r_37[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_86 = result_reg_r_37[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_87 = result_reg_r_37[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_88 = result_reg_r_37[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_89 = result_reg_r_37[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_90 = result_reg_r_37[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_91 = result_reg_r_37[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_92 = result_reg_r_37[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_93 = result_reg_r_37[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_94 = result_reg_r_37[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_95 = result_reg_r_37[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_96 = result_reg_r_37[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_97 = result_reg_r_37[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_98 = result_reg_r_37[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_99 = result_reg_r_37[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_100 = result_reg_r_37[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_101 = result_reg_r_37[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_102 = result_reg_r_37[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_103 = result_reg_r_37[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_104 = result_reg_r_37[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_75_105 = result_reg_r_37[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_38_hi_hi_hi_lo = {wire_res_75_98,wire_res_75_97,wire_res_75_96,wire_res_75_95,wire_res_75_94,
    wire_res_75_93,wire_res_75_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_38_hi_hi_lo_lo = {wire_res_75_84,wire_res_75_83,wire_res_75_82,wire_res_75_81,wire_res_75_80,
    wire_res_75_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_38_hi_hi_lo = {wire_res_75_91,wire_res_75_90,wire_res_75_89,wire_res_75_88,wire_res_75_87,
    wire_res_75_86,wire_res_75_85,result_reg_w_38_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_38_hi_lo_hi_lo = {wire_res_75_71,wire_res_75_70,wire_res_75_69,wire_res_75_68,wire_res_75_67,
    wire_res_75_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_38_hi_lo_lo_lo = {wire_res_75_58,wire_res_75_57,wire_res_75_56,wire_res_75_55,wire_res_75_54,
    wire_res_75_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_38_hi_lo_lo = {wire_res_75_65,wire_res_75_64,wire_res_75_63,wire_res_75_62,wire_res_75_61,
    wire_res_75_60,wire_res_75_59,result_reg_w_38_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_38_hi_lo = {wire_res_75_78,wire_res_75_77,wire_res_75_76,wire_res_75_75,wire_res_75_74,
    wire_res_75_73,wire_res_75_72,result_reg_w_38_hi_lo_hi_lo,result_reg_w_38_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_38_hi = {wire_res_75_105,wire_res_75_104,wire_res_75_103,wire_res_75_102,wire_res_75_101,
    wire_res_75_100,wire_res_75_99,result_reg_w_38_hi_hi_hi_lo,result_reg_w_38_hi_hi_lo,result_reg_w_38_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_38_lo_hi_hi_lo = {wire_res_75_45,wire_res_75_44,wire_res_75_43,wire_res_75_42,wire_res_75_41,
    wire_res_75_40,wire_res_75_39}; // @[BinaryDesigns2.scala 231:46]
  wire [134:0] _T_11388 = {b_aux_reg_r_37, 29'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [134:0] _GEN_1309 = {{29'd0}, a_aux_reg_r_37}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_75_29 = _GEN_1309 >= _T_11388; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_38_lo_hi_lo_lo = {wire_res_75_31,wire_res_75_30,wire_res_75_29,wire_res_75_28,wire_res_75_27,
    wire_res_75_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_38_lo_hi_lo = {wire_res_75_38,wire_res_75_37,wire_res_75_36,wire_res_75_35,wire_res_75_34,
    wire_res_75_33,wire_res_75_32,result_reg_w_38_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_38_lo_lo_hi_lo = {wire_res_75_18,wire_res_75_17,wire_res_75_16,wire_res_75_15,wire_res_75_14,
    wire_res_75_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_38_lo_lo_lo_lo = {wire_res_75_5,wire_res_75_4,wire_res_75_3,wire_res_75_2,wire_res_75_1,
    wire_res_75_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_38_lo_lo_lo = {wire_res_75_12,wire_res_75_11,wire_res_75_10,wire_res_75_9,wire_res_75_8,
    wire_res_75_7,wire_res_75_6,result_reg_w_38_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_38_lo_lo = {wire_res_75_25,wire_res_75_24,wire_res_75_23,wire_res_75_22,wire_res_75_21,
    wire_res_75_20,wire_res_75_19,result_reg_w_38_lo_lo_hi_lo,result_reg_w_38_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_38_lo = {wire_res_75_52,wire_res_75_51,wire_res_75_50,wire_res_75_49,wire_res_75_48,
    wire_res_75_47,wire_res_75_46,result_reg_w_38_lo_hi_hi_lo,result_reg_w_38_lo_hi_lo,result_reg_w_38_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_38 = {result_reg_w_38_hi,result_reg_w_38_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_76_0 = result_reg_w_38[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_1 = result_reg_w_38[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_2 = result_reg_w_38[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_3 = result_reg_w_38[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_4 = result_reg_w_38[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_5 = result_reg_w_38[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_6 = result_reg_w_38[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_7 = result_reg_w_38[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_8 = result_reg_w_38[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_9 = result_reg_w_38[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_10 = result_reg_w_38[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_11 = result_reg_w_38[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_12 = result_reg_w_38[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_13 = result_reg_w_38[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_14 = result_reg_w_38[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_15 = result_reg_w_38[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_16 = result_reg_w_38[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_17 = result_reg_w_38[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_18 = result_reg_w_38[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_19 = result_reg_w_38[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_20 = result_reg_w_38[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_21 = result_reg_w_38[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_22 = result_reg_w_38[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_23 = result_reg_w_38[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_24 = result_reg_w_38[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_25 = result_reg_w_38[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_26 = result_reg_w_38[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_27 = result_reg_w_38[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_29 = result_reg_w_38[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_30 = result_reg_w_38[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_31 = result_reg_w_38[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_32 = result_reg_w_38[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_33 = result_reg_w_38[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_34 = result_reg_w_38[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_35 = result_reg_w_38[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_36 = result_reg_w_38[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_37 = result_reg_w_38[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_38 = result_reg_w_38[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_39 = result_reg_w_38[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_40 = result_reg_w_38[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_41 = result_reg_w_38[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_42 = result_reg_w_38[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_43 = result_reg_w_38[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_44 = result_reg_w_38[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_45 = result_reg_w_38[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_46 = result_reg_w_38[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_47 = result_reg_w_38[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_48 = result_reg_w_38[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_49 = result_reg_w_38[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_50 = result_reg_w_38[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_51 = result_reg_w_38[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_52 = result_reg_w_38[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_53 = result_reg_w_38[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_54 = result_reg_w_38[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_55 = result_reg_w_38[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_56 = result_reg_w_38[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_57 = result_reg_w_38[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_58 = result_reg_w_38[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_59 = result_reg_w_38[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_60 = result_reg_w_38[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_61 = result_reg_w_38[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_62 = result_reg_w_38[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_63 = result_reg_w_38[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_64 = result_reg_w_38[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_65 = result_reg_w_38[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_66 = result_reg_w_38[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_67 = result_reg_w_38[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_68 = result_reg_w_38[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_69 = result_reg_w_38[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_70 = result_reg_w_38[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_71 = result_reg_w_38[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_72 = result_reg_w_38[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_73 = result_reg_w_38[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_74 = result_reg_w_38[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_75 = result_reg_w_38[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_76 = result_reg_w_38[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_77 = result_reg_w_38[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_78 = result_reg_w_38[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_79 = result_reg_w_38[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_80 = result_reg_w_38[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_81 = result_reg_w_38[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_82 = result_reg_w_38[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_83 = result_reg_w_38[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_84 = result_reg_w_38[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_85 = result_reg_w_38[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_86 = result_reg_w_38[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_87 = result_reg_w_38[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_88 = result_reg_w_38[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_89 = result_reg_w_38[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_90 = result_reg_w_38[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_91 = result_reg_w_38[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_92 = result_reg_w_38[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_93 = result_reg_w_38[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_94 = result_reg_w_38[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_95 = result_reg_w_38[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_96 = result_reg_w_38[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_97 = result_reg_w_38[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_98 = result_reg_w_38[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_99 = result_reg_w_38[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_100 = result_reg_w_38[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_101 = result_reg_w_38[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_102 = result_reg_w_38[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_103 = result_reg_w_38[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_104 = result_reg_w_38[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_76_105 = result_reg_w_38[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_0 = result_reg_r_38[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_1 = result_reg_r_38[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_2 = result_reg_r_38[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_3 = result_reg_r_38[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_4 = result_reg_r_38[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_5 = result_reg_r_38[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_6 = result_reg_r_38[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_7 = result_reg_r_38[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_8 = result_reg_r_38[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_9 = result_reg_r_38[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_10 = result_reg_r_38[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_11 = result_reg_r_38[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_12 = result_reg_r_38[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_13 = result_reg_r_38[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_14 = result_reg_r_38[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_15 = result_reg_r_38[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_16 = result_reg_r_38[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_17 = result_reg_r_38[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_18 = result_reg_r_38[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_19 = result_reg_r_38[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_20 = result_reg_r_38[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_21 = result_reg_r_38[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_22 = result_reg_r_38[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_23 = result_reg_r_38[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_24 = result_reg_r_38[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_25 = result_reg_r_38[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_26 = result_reg_r_38[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_28 = result_reg_r_38[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_29 = result_reg_r_38[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_30 = result_reg_r_38[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_31 = result_reg_r_38[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_32 = result_reg_r_38[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_33 = result_reg_r_38[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_34 = result_reg_r_38[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_35 = result_reg_r_38[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_36 = result_reg_r_38[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_37 = result_reg_r_38[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_38 = result_reg_r_38[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_39 = result_reg_r_38[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_40 = result_reg_r_38[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_41 = result_reg_r_38[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_42 = result_reg_r_38[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_43 = result_reg_r_38[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_44 = result_reg_r_38[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_45 = result_reg_r_38[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_46 = result_reg_r_38[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_47 = result_reg_r_38[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_48 = result_reg_r_38[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_49 = result_reg_r_38[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_50 = result_reg_r_38[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_51 = result_reg_r_38[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_52 = result_reg_r_38[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_53 = result_reg_r_38[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_54 = result_reg_r_38[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_55 = result_reg_r_38[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_56 = result_reg_r_38[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_57 = result_reg_r_38[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_58 = result_reg_r_38[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_59 = result_reg_r_38[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_60 = result_reg_r_38[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_61 = result_reg_r_38[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_62 = result_reg_r_38[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_63 = result_reg_r_38[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_64 = result_reg_r_38[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_65 = result_reg_r_38[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_66 = result_reg_r_38[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_67 = result_reg_r_38[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_68 = result_reg_r_38[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_69 = result_reg_r_38[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_70 = result_reg_r_38[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_71 = result_reg_r_38[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_72 = result_reg_r_38[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_73 = result_reg_r_38[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_74 = result_reg_r_38[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_75 = result_reg_r_38[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_76 = result_reg_r_38[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_77 = result_reg_r_38[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_78 = result_reg_r_38[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_79 = result_reg_r_38[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_80 = result_reg_r_38[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_81 = result_reg_r_38[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_82 = result_reg_r_38[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_83 = result_reg_r_38[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_84 = result_reg_r_38[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_85 = result_reg_r_38[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_86 = result_reg_r_38[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_87 = result_reg_r_38[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_88 = result_reg_r_38[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_89 = result_reg_r_38[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_90 = result_reg_r_38[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_91 = result_reg_r_38[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_92 = result_reg_r_38[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_93 = result_reg_r_38[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_94 = result_reg_r_38[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_95 = result_reg_r_38[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_96 = result_reg_r_38[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_97 = result_reg_r_38[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_98 = result_reg_r_38[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_99 = result_reg_r_38[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_100 = result_reg_r_38[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_101 = result_reg_r_38[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_102 = result_reg_r_38[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_103 = result_reg_r_38[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_104 = result_reg_r_38[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_77_105 = result_reg_r_38[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_39_hi_hi_hi_lo = {wire_res_77_98,wire_res_77_97,wire_res_77_96,wire_res_77_95,wire_res_77_94,
    wire_res_77_93,wire_res_77_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_39_hi_hi_lo_lo = {wire_res_77_84,wire_res_77_83,wire_res_77_82,wire_res_77_81,wire_res_77_80,
    wire_res_77_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_39_hi_hi_lo = {wire_res_77_91,wire_res_77_90,wire_res_77_89,wire_res_77_88,wire_res_77_87,
    wire_res_77_86,wire_res_77_85,result_reg_w_39_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_39_hi_lo_hi_lo = {wire_res_77_71,wire_res_77_70,wire_res_77_69,wire_res_77_68,wire_res_77_67,
    wire_res_77_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_39_hi_lo_lo_lo = {wire_res_77_58,wire_res_77_57,wire_res_77_56,wire_res_77_55,wire_res_77_54,
    wire_res_77_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_39_hi_lo_lo = {wire_res_77_65,wire_res_77_64,wire_res_77_63,wire_res_77_62,wire_res_77_61,
    wire_res_77_60,wire_res_77_59,result_reg_w_39_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_39_hi_lo = {wire_res_77_78,wire_res_77_77,wire_res_77_76,wire_res_77_75,wire_res_77_74,
    wire_res_77_73,wire_res_77_72,result_reg_w_39_hi_lo_hi_lo,result_reg_w_39_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_39_hi = {wire_res_77_105,wire_res_77_104,wire_res_77_103,wire_res_77_102,wire_res_77_101,
    wire_res_77_100,wire_res_77_99,result_reg_w_39_hi_hi_hi_lo,result_reg_w_39_hi_hi_lo,result_reg_w_39_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_39_lo_hi_hi_lo = {wire_res_77_45,wire_res_77_44,wire_res_77_43,wire_res_77_42,wire_res_77_41,
    wire_res_77_40,wire_res_77_39}; // @[BinaryDesigns2.scala 231:46]
  wire [132:0] _T_11392 = {b_aux_reg_r_38, 27'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [132:0] _GEN_1310 = {{27'd0}, a_aux_reg_r_38}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_77_27 = _GEN_1310 >= _T_11392; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_39_lo_hi_lo_lo = {wire_res_77_31,wire_res_77_30,wire_res_77_29,wire_res_77_28,wire_res_77_27,
    wire_res_77_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_39_lo_hi_lo = {wire_res_77_38,wire_res_77_37,wire_res_77_36,wire_res_77_35,wire_res_77_34,
    wire_res_77_33,wire_res_77_32,result_reg_w_39_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_39_lo_lo_hi_lo = {wire_res_77_18,wire_res_77_17,wire_res_77_16,wire_res_77_15,wire_res_77_14,
    wire_res_77_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_39_lo_lo_lo_lo = {wire_res_77_5,wire_res_77_4,wire_res_77_3,wire_res_77_2,wire_res_77_1,
    wire_res_77_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_39_lo_lo_lo = {wire_res_77_12,wire_res_77_11,wire_res_77_10,wire_res_77_9,wire_res_77_8,
    wire_res_77_7,wire_res_77_6,result_reg_w_39_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_39_lo_lo = {wire_res_77_25,wire_res_77_24,wire_res_77_23,wire_res_77_22,wire_res_77_21,
    wire_res_77_20,wire_res_77_19,result_reg_w_39_lo_lo_hi_lo,result_reg_w_39_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_39_lo = {wire_res_77_52,wire_res_77_51,wire_res_77_50,wire_res_77_49,wire_res_77_48,
    wire_res_77_47,wire_res_77_46,result_reg_w_39_lo_hi_hi_lo,result_reg_w_39_lo_hi_lo,result_reg_w_39_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_39 = {result_reg_w_39_hi,result_reg_w_39_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_78_0 = result_reg_w_39[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_1 = result_reg_w_39[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_2 = result_reg_w_39[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_3 = result_reg_w_39[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_4 = result_reg_w_39[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_5 = result_reg_w_39[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_6 = result_reg_w_39[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_7 = result_reg_w_39[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_8 = result_reg_w_39[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_9 = result_reg_w_39[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_10 = result_reg_w_39[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_11 = result_reg_w_39[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_12 = result_reg_w_39[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_13 = result_reg_w_39[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_14 = result_reg_w_39[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_15 = result_reg_w_39[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_16 = result_reg_w_39[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_17 = result_reg_w_39[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_18 = result_reg_w_39[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_19 = result_reg_w_39[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_20 = result_reg_w_39[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_21 = result_reg_w_39[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_22 = result_reg_w_39[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_23 = result_reg_w_39[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_24 = result_reg_w_39[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_25 = result_reg_w_39[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_27 = result_reg_w_39[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_28 = result_reg_w_39[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_29 = result_reg_w_39[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_30 = result_reg_w_39[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_31 = result_reg_w_39[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_32 = result_reg_w_39[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_33 = result_reg_w_39[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_34 = result_reg_w_39[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_35 = result_reg_w_39[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_36 = result_reg_w_39[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_37 = result_reg_w_39[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_38 = result_reg_w_39[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_39 = result_reg_w_39[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_40 = result_reg_w_39[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_41 = result_reg_w_39[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_42 = result_reg_w_39[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_43 = result_reg_w_39[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_44 = result_reg_w_39[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_45 = result_reg_w_39[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_46 = result_reg_w_39[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_47 = result_reg_w_39[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_48 = result_reg_w_39[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_49 = result_reg_w_39[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_50 = result_reg_w_39[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_51 = result_reg_w_39[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_52 = result_reg_w_39[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_53 = result_reg_w_39[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_54 = result_reg_w_39[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_55 = result_reg_w_39[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_56 = result_reg_w_39[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_57 = result_reg_w_39[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_58 = result_reg_w_39[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_59 = result_reg_w_39[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_60 = result_reg_w_39[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_61 = result_reg_w_39[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_62 = result_reg_w_39[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_63 = result_reg_w_39[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_64 = result_reg_w_39[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_65 = result_reg_w_39[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_66 = result_reg_w_39[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_67 = result_reg_w_39[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_68 = result_reg_w_39[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_69 = result_reg_w_39[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_70 = result_reg_w_39[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_71 = result_reg_w_39[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_72 = result_reg_w_39[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_73 = result_reg_w_39[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_74 = result_reg_w_39[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_75 = result_reg_w_39[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_76 = result_reg_w_39[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_77 = result_reg_w_39[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_78 = result_reg_w_39[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_79 = result_reg_w_39[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_80 = result_reg_w_39[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_81 = result_reg_w_39[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_82 = result_reg_w_39[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_83 = result_reg_w_39[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_84 = result_reg_w_39[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_85 = result_reg_w_39[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_86 = result_reg_w_39[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_87 = result_reg_w_39[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_88 = result_reg_w_39[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_89 = result_reg_w_39[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_90 = result_reg_w_39[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_91 = result_reg_w_39[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_92 = result_reg_w_39[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_93 = result_reg_w_39[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_94 = result_reg_w_39[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_95 = result_reg_w_39[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_96 = result_reg_w_39[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_97 = result_reg_w_39[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_98 = result_reg_w_39[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_99 = result_reg_w_39[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_100 = result_reg_w_39[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_101 = result_reg_w_39[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_102 = result_reg_w_39[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_103 = result_reg_w_39[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_104 = result_reg_w_39[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_78_105 = result_reg_w_39[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_0 = result_reg_r_39[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_1 = result_reg_r_39[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_2 = result_reg_r_39[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_3 = result_reg_r_39[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_4 = result_reg_r_39[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_5 = result_reg_r_39[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_6 = result_reg_r_39[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_7 = result_reg_r_39[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_8 = result_reg_r_39[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_9 = result_reg_r_39[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_10 = result_reg_r_39[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_11 = result_reg_r_39[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_12 = result_reg_r_39[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_13 = result_reg_r_39[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_14 = result_reg_r_39[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_15 = result_reg_r_39[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_16 = result_reg_r_39[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_17 = result_reg_r_39[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_18 = result_reg_r_39[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_19 = result_reg_r_39[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_20 = result_reg_r_39[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_21 = result_reg_r_39[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_22 = result_reg_r_39[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_23 = result_reg_r_39[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_24 = result_reg_r_39[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_26 = result_reg_r_39[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_27 = result_reg_r_39[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_28 = result_reg_r_39[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_29 = result_reg_r_39[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_30 = result_reg_r_39[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_31 = result_reg_r_39[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_32 = result_reg_r_39[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_33 = result_reg_r_39[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_34 = result_reg_r_39[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_35 = result_reg_r_39[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_36 = result_reg_r_39[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_37 = result_reg_r_39[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_38 = result_reg_r_39[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_39 = result_reg_r_39[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_40 = result_reg_r_39[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_41 = result_reg_r_39[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_42 = result_reg_r_39[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_43 = result_reg_r_39[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_44 = result_reg_r_39[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_45 = result_reg_r_39[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_46 = result_reg_r_39[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_47 = result_reg_r_39[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_48 = result_reg_r_39[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_49 = result_reg_r_39[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_50 = result_reg_r_39[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_51 = result_reg_r_39[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_52 = result_reg_r_39[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_53 = result_reg_r_39[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_54 = result_reg_r_39[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_55 = result_reg_r_39[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_56 = result_reg_r_39[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_57 = result_reg_r_39[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_58 = result_reg_r_39[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_59 = result_reg_r_39[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_60 = result_reg_r_39[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_61 = result_reg_r_39[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_62 = result_reg_r_39[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_63 = result_reg_r_39[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_64 = result_reg_r_39[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_65 = result_reg_r_39[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_66 = result_reg_r_39[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_67 = result_reg_r_39[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_68 = result_reg_r_39[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_69 = result_reg_r_39[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_70 = result_reg_r_39[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_71 = result_reg_r_39[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_72 = result_reg_r_39[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_73 = result_reg_r_39[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_74 = result_reg_r_39[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_75 = result_reg_r_39[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_76 = result_reg_r_39[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_77 = result_reg_r_39[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_78 = result_reg_r_39[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_79 = result_reg_r_39[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_80 = result_reg_r_39[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_81 = result_reg_r_39[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_82 = result_reg_r_39[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_83 = result_reg_r_39[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_84 = result_reg_r_39[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_85 = result_reg_r_39[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_86 = result_reg_r_39[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_87 = result_reg_r_39[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_88 = result_reg_r_39[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_89 = result_reg_r_39[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_90 = result_reg_r_39[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_91 = result_reg_r_39[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_92 = result_reg_r_39[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_93 = result_reg_r_39[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_94 = result_reg_r_39[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_95 = result_reg_r_39[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_96 = result_reg_r_39[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_97 = result_reg_r_39[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_98 = result_reg_r_39[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_99 = result_reg_r_39[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_100 = result_reg_r_39[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_101 = result_reg_r_39[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_102 = result_reg_r_39[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_103 = result_reg_r_39[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_104 = result_reg_r_39[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_79_105 = result_reg_r_39[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_40_hi_hi_hi_lo = {wire_res_79_98,wire_res_79_97,wire_res_79_96,wire_res_79_95,wire_res_79_94,
    wire_res_79_93,wire_res_79_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_40_hi_hi_lo_lo = {wire_res_79_84,wire_res_79_83,wire_res_79_82,wire_res_79_81,wire_res_79_80,
    wire_res_79_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_40_hi_hi_lo = {wire_res_79_91,wire_res_79_90,wire_res_79_89,wire_res_79_88,wire_res_79_87,
    wire_res_79_86,wire_res_79_85,result_reg_w_40_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_40_hi_lo_hi_lo = {wire_res_79_71,wire_res_79_70,wire_res_79_69,wire_res_79_68,wire_res_79_67,
    wire_res_79_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_40_hi_lo_lo_lo = {wire_res_79_58,wire_res_79_57,wire_res_79_56,wire_res_79_55,wire_res_79_54,
    wire_res_79_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_40_hi_lo_lo = {wire_res_79_65,wire_res_79_64,wire_res_79_63,wire_res_79_62,wire_res_79_61,
    wire_res_79_60,wire_res_79_59,result_reg_w_40_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_40_hi_lo = {wire_res_79_78,wire_res_79_77,wire_res_79_76,wire_res_79_75,wire_res_79_74,
    wire_res_79_73,wire_res_79_72,result_reg_w_40_hi_lo_hi_lo,result_reg_w_40_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_40_hi = {wire_res_79_105,wire_res_79_104,wire_res_79_103,wire_res_79_102,wire_res_79_101,
    wire_res_79_100,wire_res_79_99,result_reg_w_40_hi_hi_hi_lo,result_reg_w_40_hi_hi_lo,result_reg_w_40_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_40_lo_hi_hi_lo = {wire_res_79_45,wire_res_79_44,wire_res_79_43,wire_res_79_42,wire_res_79_41,
    wire_res_79_40,wire_res_79_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_40_lo_hi_lo_lo = {wire_res_79_31,wire_res_79_30,wire_res_79_29,wire_res_79_28,wire_res_79_27,
    wire_res_79_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_40_lo_hi_lo = {wire_res_79_38,wire_res_79_37,wire_res_79_36,wire_res_79_35,wire_res_79_34,
    wire_res_79_33,wire_res_79_32,result_reg_w_40_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [130:0] _T_11396 = {b_aux_reg_r_39, 25'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [130:0] _GEN_1311 = {{25'd0}, a_aux_reg_r_39}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_79_25 = _GEN_1311 >= _T_11396; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_40_lo_lo_hi_lo = {wire_res_79_18,wire_res_79_17,wire_res_79_16,wire_res_79_15,wire_res_79_14,
    wire_res_79_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_40_lo_lo_lo_lo = {wire_res_79_5,wire_res_79_4,wire_res_79_3,wire_res_79_2,wire_res_79_1,
    wire_res_79_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_40_lo_lo_lo = {wire_res_79_12,wire_res_79_11,wire_res_79_10,wire_res_79_9,wire_res_79_8,
    wire_res_79_7,wire_res_79_6,result_reg_w_40_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_40_lo_lo = {wire_res_79_25,wire_res_79_24,wire_res_79_23,wire_res_79_22,wire_res_79_21,
    wire_res_79_20,wire_res_79_19,result_reg_w_40_lo_lo_hi_lo,result_reg_w_40_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_40_lo = {wire_res_79_52,wire_res_79_51,wire_res_79_50,wire_res_79_49,wire_res_79_48,
    wire_res_79_47,wire_res_79_46,result_reg_w_40_lo_hi_hi_lo,result_reg_w_40_lo_hi_lo,result_reg_w_40_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_40 = {result_reg_w_40_hi,result_reg_w_40_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_80_0 = result_reg_w_40[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_1 = result_reg_w_40[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_2 = result_reg_w_40[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_3 = result_reg_w_40[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_4 = result_reg_w_40[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_5 = result_reg_w_40[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_6 = result_reg_w_40[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_7 = result_reg_w_40[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_8 = result_reg_w_40[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_9 = result_reg_w_40[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_10 = result_reg_w_40[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_11 = result_reg_w_40[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_12 = result_reg_w_40[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_13 = result_reg_w_40[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_14 = result_reg_w_40[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_15 = result_reg_w_40[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_16 = result_reg_w_40[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_17 = result_reg_w_40[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_18 = result_reg_w_40[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_19 = result_reg_w_40[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_20 = result_reg_w_40[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_21 = result_reg_w_40[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_22 = result_reg_w_40[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_23 = result_reg_w_40[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_25 = result_reg_w_40[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_26 = result_reg_w_40[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_27 = result_reg_w_40[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_28 = result_reg_w_40[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_29 = result_reg_w_40[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_30 = result_reg_w_40[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_31 = result_reg_w_40[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_32 = result_reg_w_40[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_33 = result_reg_w_40[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_34 = result_reg_w_40[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_35 = result_reg_w_40[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_36 = result_reg_w_40[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_37 = result_reg_w_40[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_38 = result_reg_w_40[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_39 = result_reg_w_40[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_40 = result_reg_w_40[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_41 = result_reg_w_40[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_42 = result_reg_w_40[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_43 = result_reg_w_40[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_44 = result_reg_w_40[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_45 = result_reg_w_40[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_46 = result_reg_w_40[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_47 = result_reg_w_40[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_48 = result_reg_w_40[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_49 = result_reg_w_40[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_50 = result_reg_w_40[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_51 = result_reg_w_40[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_52 = result_reg_w_40[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_53 = result_reg_w_40[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_54 = result_reg_w_40[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_55 = result_reg_w_40[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_56 = result_reg_w_40[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_57 = result_reg_w_40[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_58 = result_reg_w_40[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_59 = result_reg_w_40[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_60 = result_reg_w_40[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_61 = result_reg_w_40[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_62 = result_reg_w_40[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_63 = result_reg_w_40[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_64 = result_reg_w_40[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_65 = result_reg_w_40[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_66 = result_reg_w_40[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_67 = result_reg_w_40[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_68 = result_reg_w_40[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_69 = result_reg_w_40[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_70 = result_reg_w_40[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_71 = result_reg_w_40[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_72 = result_reg_w_40[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_73 = result_reg_w_40[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_74 = result_reg_w_40[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_75 = result_reg_w_40[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_76 = result_reg_w_40[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_77 = result_reg_w_40[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_78 = result_reg_w_40[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_79 = result_reg_w_40[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_80 = result_reg_w_40[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_81 = result_reg_w_40[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_82 = result_reg_w_40[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_83 = result_reg_w_40[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_84 = result_reg_w_40[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_85 = result_reg_w_40[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_86 = result_reg_w_40[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_87 = result_reg_w_40[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_88 = result_reg_w_40[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_89 = result_reg_w_40[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_90 = result_reg_w_40[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_91 = result_reg_w_40[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_92 = result_reg_w_40[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_93 = result_reg_w_40[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_94 = result_reg_w_40[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_95 = result_reg_w_40[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_96 = result_reg_w_40[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_97 = result_reg_w_40[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_98 = result_reg_w_40[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_99 = result_reg_w_40[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_100 = result_reg_w_40[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_101 = result_reg_w_40[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_102 = result_reg_w_40[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_103 = result_reg_w_40[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_104 = result_reg_w_40[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_80_105 = result_reg_w_40[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_0 = result_reg_r_40[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_1 = result_reg_r_40[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_2 = result_reg_r_40[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_3 = result_reg_r_40[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_4 = result_reg_r_40[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_5 = result_reg_r_40[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_6 = result_reg_r_40[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_7 = result_reg_r_40[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_8 = result_reg_r_40[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_9 = result_reg_r_40[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_10 = result_reg_r_40[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_11 = result_reg_r_40[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_12 = result_reg_r_40[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_13 = result_reg_r_40[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_14 = result_reg_r_40[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_15 = result_reg_r_40[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_16 = result_reg_r_40[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_17 = result_reg_r_40[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_18 = result_reg_r_40[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_19 = result_reg_r_40[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_20 = result_reg_r_40[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_21 = result_reg_r_40[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_22 = result_reg_r_40[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_24 = result_reg_r_40[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_25 = result_reg_r_40[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_26 = result_reg_r_40[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_27 = result_reg_r_40[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_28 = result_reg_r_40[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_29 = result_reg_r_40[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_30 = result_reg_r_40[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_31 = result_reg_r_40[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_32 = result_reg_r_40[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_33 = result_reg_r_40[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_34 = result_reg_r_40[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_35 = result_reg_r_40[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_36 = result_reg_r_40[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_37 = result_reg_r_40[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_38 = result_reg_r_40[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_39 = result_reg_r_40[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_40 = result_reg_r_40[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_41 = result_reg_r_40[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_42 = result_reg_r_40[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_43 = result_reg_r_40[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_44 = result_reg_r_40[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_45 = result_reg_r_40[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_46 = result_reg_r_40[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_47 = result_reg_r_40[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_48 = result_reg_r_40[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_49 = result_reg_r_40[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_50 = result_reg_r_40[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_51 = result_reg_r_40[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_52 = result_reg_r_40[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_53 = result_reg_r_40[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_54 = result_reg_r_40[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_55 = result_reg_r_40[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_56 = result_reg_r_40[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_57 = result_reg_r_40[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_58 = result_reg_r_40[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_59 = result_reg_r_40[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_60 = result_reg_r_40[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_61 = result_reg_r_40[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_62 = result_reg_r_40[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_63 = result_reg_r_40[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_64 = result_reg_r_40[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_65 = result_reg_r_40[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_66 = result_reg_r_40[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_67 = result_reg_r_40[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_68 = result_reg_r_40[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_69 = result_reg_r_40[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_70 = result_reg_r_40[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_71 = result_reg_r_40[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_72 = result_reg_r_40[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_73 = result_reg_r_40[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_74 = result_reg_r_40[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_75 = result_reg_r_40[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_76 = result_reg_r_40[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_77 = result_reg_r_40[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_78 = result_reg_r_40[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_79 = result_reg_r_40[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_80 = result_reg_r_40[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_81 = result_reg_r_40[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_82 = result_reg_r_40[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_83 = result_reg_r_40[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_84 = result_reg_r_40[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_85 = result_reg_r_40[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_86 = result_reg_r_40[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_87 = result_reg_r_40[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_88 = result_reg_r_40[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_89 = result_reg_r_40[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_90 = result_reg_r_40[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_91 = result_reg_r_40[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_92 = result_reg_r_40[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_93 = result_reg_r_40[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_94 = result_reg_r_40[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_95 = result_reg_r_40[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_96 = result_reg_r_40[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_97 = result_reg_r_40[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_98 = result_reg_r_40[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_99 = result_reg_r_40[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_100 = result_reg_r_40[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_101 = result_reg_r_40[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_102 = result_reg_r_40[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_103 = result_reg_r_40[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_104 = result_reg_r_40[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_81_105 = result_reg_r_40[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_41_hi_hi_hi_lo = {wire_res_81_98,wire_res_81_97,wire_res_81_96,wire_res_81_95,wire_res_81_94,
    wire_res_81_93,wire_res_81_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_41_hi_hi_lo_lo = {wire_res_81_84,wire_res_81_83,wire_res_81_82,wire_res_81_81,wire_res_81_80,
    wire_res_81_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_41_hi_hi_lo = {wire_res_81_91,wire_res_81_90,wire_res_81_89,wire_res_81_88,wire_res_81_87,
    wire_res_81_86,wire_res_81_85,result_reg_w_41_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_41_hi_lo_hi_lo = {wire_res_81_71,wire_res_81_70,wire_res_81_69,wire_res_81_68,wire_res_81_67,
    wire_res_81_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_41_hi_lo_lo_lo = {wire_res_81_58,wire_res_81_57,wire_res_81_56,wire_res_81_55,wire_res_81_54,
    wire_res_81_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_41_hi_lo_lo = {wire_res_81_65,wire_res_81_64,wire_res_81_63,wire_res_81_62,wire_res_81_61,
    wire_res_81_60,wire_res_81_59,result_reg_w_41_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_41_hi_lo = {wire_res_81_78,wire_res_81_77,wire_res_81_76,wire_res_81_75,wire_res_81_74,
    wire_res_81_73,wire_res_81_72,result_reg_w_41_hi_lo_hi_lo,result_reg_w_41_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_41_hi = {wire_res_81_105,wire_res_81_104,wire_res_81_103,wire_res_81_102,wire_res_81_101,
    wire_res_81_100,wire_res_81_99,result_reg_w_41_hi_hi_hi_lo,result_reg_w_41_hi_hi_lo,result_reg_w_41_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_41_lo_hi_hi_lo = {wire_res_81_45,wire_res_81_44,wire_res_81_43,wire_res_81_42,wire_res_81_41,
    wire_res_81_40,wire_res_81_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_41_lo_hi_lo_lo = {wire_res_81_31,wire_res_81_30,wire_res_81_29,wire_res_81_28,wire_res_81_27,
    wire_res_81_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_41_lo_hi_lo = {wire_res_81_38,wire_res_81_37,wire_res_81_36,wire_res_81_35,wire_res_81_34,
    wire_res_81_33,wire_res_81_32,result_reg_w_41_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [128:0] _T_11400 = {b_aux_reg_r_40, 23'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [128:0] _GEN_1312 = {{23'd0}, a_aux_reg_r_40}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_81_23 = _GEN_1312 >= _T_11400; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_41_lo_lo_hi_lo = {wire_res_81_18,wire_res_81_17,wire_res_81_16,wire_res_81_15,wire_res_81_14,
    wire_res_81_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_41_lo_lo_lo_lo = {wire_res_81_5,wire_res_81_4,wire_res_81_3,wire_res_81_2,wire_res_81_1,
    wire_res_81_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_41_lo_lo_lo = {wire_res_81_12,wire_res_81_11,wire_res_81_10,wire_res_81_9,wire_res_81_8,
    wire_res_81_7,wire_res_81_6,result_reg_w_41_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_41_lo_lo = {wire_res_81_25,wire_res_81_24,wire_res_81_23,wire_res_81_22,wire_res_81_21,
    wire_res_81_20,wire_res_81_19,result_reg_w_41_lo_lo_hi_lo,result_reg_w_41_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_41_lo = {wire_res_81_52,wire_res_81_51,wire_res_81_50,wire_res_81_49,wire_res_81_48,
    wire_res_81_47,wire_res_81_46,result_reg_w_41_lo_hi_hi_lo,result_reg_w_41_lo_hi_lo,result_reg_w_41_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_41 = {result_reg_w_41_hi,result_reg_w_41_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_82_0 = result_reg_w_41[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_1 = result_reg_w_41[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_2 = result_reg_w_41[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_3 = result_reg_w_41[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_4 = result_reg_w_41[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_5 = result_reg_w_41[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_6 = result_reg_w_41[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_7 = result_reg_w_41[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_8 = result_reg_w_41[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_9 = result_reg_w_41[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_10 = result_reg_w_41[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_11 = result_reg_w_41[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_12 = result_reg_w_41[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_13 = result_reg_w_41[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_14 = result_reg_w_41[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_15 = result_reg_w_41[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_16 = result_reg_w_41[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_17 = result_reg_w_41[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_18 = result_reg_w_41[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_19 = result_reg_w_41[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_20 = result_reg_w_41[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_21 = result_reg_w_41[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_23 = result_reg_w_41[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_24 = result_reg_w_41[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_25 = result_reg_w_41[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_26 = result_reg_w_41[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_27 = result_reg_w_41[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_28 = result_reg_w_41[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_29 = result_reg_w_41[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_30 = result_reg_w_41[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_31 = result_reg_w_41[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_32 = result_reg_w_41[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_33 = result_reg_w_41[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_34 = result_reg_w_41[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_35 = result_reg_w_41[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_36 = result_reg_w_41[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_37 = result_reg_w_41[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_38 = result_reg_w_41[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_39 = result_reg_w_41[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_40 = result_reg_w_41[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_41 = result_reg_w_41[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_42 = result_reg_w_41[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_43 = result_reg_w_41[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_44 = result_reg_w_41[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_45 = result_reg_w_41[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_46 = result_reg_w_41[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_47 = result_reg_w_41[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_48 = result_reg_w_41[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_49 = result_reg_w_41[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_50 = result_reg_w_41[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_51 = result_reg_w_41[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_52 = result_reg_w_41[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_53 = result_reg_w_41[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_54 = result_reg_w_41[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_55 = result_reg_w_41[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_56 = result_reg_w_41[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_57 = result_reg_w_41[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_58 = result_reg_w_41[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_59 = result_reg_w_41[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_60 = result_reg_w_41[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_61 = result_reg_w_41[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_62 = result_reg_w_41[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_63 = result_reg_w_41[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_64 = result_reg_w_41[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_65 = result_reg_w_41[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_66 = result_reg_w_41[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_67 = result_reg_w_41[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_68 = result_reg_w_41[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_69 = result_reg_w_41[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_70 = result_reg_w_41[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_71 = result_reg_w_41[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_72 = result_reg_w_41[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_73 = result_reg_w_41[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_74 = result_reg_w_41[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_75 = result_reg_w_41[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_76 = result_reg_w_41[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_77 = result_reg_w_41[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_78 = result_reg_w_41[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_79 = result_reg_w_41[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_80 = result_reg_w_41[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_81 = result_reg_w_41[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_82 = result_reg_w_41[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_83 = result_reg_w_41[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_84 = result_reg_w_41[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_85 = result_reg_w_41[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_86 = result_reg_w_41[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_87 = result_reg_w_41[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_88 = result_reg_w_41[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_89 = result_reg_w_41[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_90 = result_reg_w_41[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_91 = result_reg_w_41[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_92 = result_reg_w_41[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_93 = result_reg_w_41[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_94 = result_reg_w_41[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_95 = result_reg_w_41[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_96 = result_reg_w_41[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_97 = result_reg_w_41[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_98 = result_reg_w_41[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_99 = result_reg_w_41[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_100 = result_reg_w_41[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_101 = result_reg_w_41[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_102 = result_reg_w_41[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_103 = result_reg_w_41[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_104 = result_reg_w_41[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_82_105 = result_reg_w_41[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_0 = result_reg_r_41[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_1 = result_reg_r_41[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_2 = result_reg_r_41[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_3 = result_reg_r_41[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_4 = result_reg_r_41[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_5 = result_reg_r_41[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_6 = result_reg_r_41[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_7 = result_reg_r_41[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_8 = result_reg_r_41[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_9 = result_reg_r_41[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_10 = result_reg_r_41[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_11 = result_reg_r_41[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_12 = result_reg_r_41[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_13 = result_reg_r_41[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_14 = result_reg_r_41[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_15 = result_reg_r_41[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_16 = result_reg_r_41[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_17 = result_reg_r_41[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_18 = result_reg_r_41[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_19 = result_reg_r_41[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_20 = result_reg_r_41[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_22 = result_reg_r_41[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_23 = result_reg_r_41[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_24 = result_reg_r_41[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_25 = result_reg_r_41[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_26 = result_reg_r_41[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_27 = result_reg_r_41[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_28 = result_reg_r_41[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_29 = result_reg_r_41[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_30 = result_reg_r_41[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_31 = result_reg_r_41[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_32 = result_reg_r_41[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_33 = result_reg_r_41[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_34 = result_reg_r_41[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_35 = result_reg_r_41[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_36 = result_reg_r_41[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_37 = result_reg_r_41[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_38 = result_reg_r_41[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_39 = result_reg_r_41[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_40 = result_reg_r_41[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_41 = result_reg_r_41[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_42 = result_reg_r_41[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_43 = result_reg_r_41[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_44 = result_reg_r_41[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_45 = result_reg_r_41[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_46 = result_reg_r_41[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_47 = result_reg_r_41[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_48 = result_reg_r_41[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_49 = result_reg_r_41[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_50 = result_reg_r_41[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_51 = result_reg_r_41[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_52 = result_reg_r_41[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_53 = result_reg_r_41[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_54 = result_reg_r_41[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_55 = result_reg_r_41[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_56 = result_reg_r_41[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_57 = result_reg_r_41[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_58 = result_reg_r_41[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_59 = result_reg_r_41[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_60 = result_reg_r_41[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_61 = result_reg_r_41[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_62 = result_reg_r_41[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_63 = result_reg_r_41[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_64 = result_reg_r_41[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_65 = result_reg_r_41[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_66 = result_reg_r_41[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_67 = result_reg_r_41[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_68 = result_reg_r_41[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_69 = result_reg_r_41[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_70 = result_reg_r_41[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_71 = result_reg_r_41[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_72 = result_reg_r_41[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_73 = result_reg_r_41[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_74 = result_reg_r_41[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_75 = result_reg_r_41[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_76 = result_reg_r_41[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_77 = result_reg_r_41[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_78 = result_reg_r_41[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_79 = result_reg_r_41[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_80 = result_reg_r_41[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_81 = result_reg_r_41[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_82 = result_reg_r_41[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_83 = result_reg_r_41[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_84 = result_reg_r_41[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_85 = result_reg_r_41[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_86 = result_reg_r_41[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_87 = result_reg_r_41[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_88 = result_reg_r_41[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_89 = result_reg_r_41[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_90 = result_reg_r_41[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_91 = result_reg_r_41[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_92 = result_reg_r_41[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_93 = result_reg_r_41[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_94 = result_reg_r_41[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_95 = result_reg_r_41[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_96 = result_reg_r_41[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_97 = result_reg_r_41[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_98 = result_reg_r_41[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_99 = result_reg_r_41[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_100 = result_reg_r_41[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_101 = result_reg_r_41[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_102 = result_reg_r_41[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_103 = result_reg_r_41[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_104 = result_reg_r_41[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_83_105 = result_reg_r_41[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_42_hi_hi_hi_lo = {wire_res_83_98,wire_res_83_97,wire_res_83_96,wire_res_83_95,wire_res_83_94,
    wire_res_83_93,wire_res_83_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_42_hi_hi_lo_lo = {wire_res_83_84,wire_res_83_83,wire_res_83_82,wire_res_83_81,wire_res_83_80,
    wire_res_83_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_42_hi_hi_lo = {wire_res_83_91,wire_res_83_90,wire_res_83_89,wire_res_83_88,wire_res_83_87,
    wire_res_83_86,wire_res_83_85,result_reg_w_42_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_42_hi_lo_hi_lo = {wire_res_83_71,wire_res_83_70,wire_res_83_69,wire_res_83_68,wire_res_83_67,
    wire_res_83_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_42_hi_lo_lo_lo = {wire_res_83_58,wire_res_83_57,wire_res_83_56,wire_res_83_55,wire_res_83_54,
    wire_res_83_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_42_hi_lo_lo = {wire_res_83_65,wire_res_83_64,wire_res_83_63,wire_res_83_62,wire_res_83_61,
    wire_res_83_60,wire_res_83_59,result_reg_w_42_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_42_hi_lo = {wire_res_83_78,wire_res_83_77,wire_res_83_76,wire_res_83_75,wire_res_83_74,
    wire_res_83_73,wire_res_83_72,result_reg_w_42_hi_lo_hi_lo,result_reg_w_42_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_42_hi = {wire_res_83_105,wire_res_83_104,wire_res_83_103,wire_res_83_102,wire_res_83_101,
    wire_res_83_100,wire_res_83_99,result_reg_w_42_hi_hi_hi_lo,result_reg_w_42_hi_hi_lo,result_reg_w_42_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_42_lo_hi_hi_lo = {wire_res_83_45,wire_res_83_44,wire_res_83_43,wire_res_83_42,wire_res_83_41,
    wire_res_83_40,wire_res_83_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_42_lo_hi_lo_lo = {wire_res_83_31,wire_res_83_30,wire_res_83_29,wire_res_83_28,wire_res_83_27,
    wire_res_83_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_42_lo_hi_lo = {wire_res_83_38,wire_res_83_37,wire_res_83_36,wire_res_83_35,wire_res_83_34,
    wire_res_83_33,wire_res_83_32,result_reg_w_42_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [126:0] _T_11404 = {b_aux_reg_r_41, 21'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [126:0] _GEN_1313 = {{21'd0}, a_aux_reg_r_41}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_83_21 = _GEN_1313 >= _T_11404; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_42_lo_lo_hi_lo = {wire_res_83_18,wire_res_83_17,wire_res_83_16,wire_res_83_15,wire_res_83_14,
    wire_res_83_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_42_lo_lo_lo_lo = {wire_res_83_5,wire_res_83_4,wire_res_83_3,wire_res_83_2,wire_res_83_1,
    wire_res_83_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_42_lo_lo_lo = {wire_res_83_12,wire_res_83_11,wire_res_83_10,wire_res_83_9,wire_res_83_8,
    wire_res_83_7,wire_res_83_6,result_reg_w_42_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_42_lo_lo = {wire_res_83_25,wire_res_83_24,wire_res_83_23,wire_res_83_22,wire_res_83_21,
    wire_res_83_20,wire_res_83_19,result_reg_w_42_lo_lo_hi_lo,result_reg_w_42_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_42_lo = {wire_res_83_52,wire_res_83_51,wire_res_83_50,wire_res_83_49,wire_res_83_48,
    wire_res_83_47,wire_res_83_46,result_reg_w_42_lo_hi_hi_lo,result_reg_w_42_lo_hi_lo,result_reg_w_42_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_42 = {result_reg_w_42_hi,result_reg_w_42_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_84_0 = result_reg_w_42[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_1 = result_reg_w_42[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_2 = result_reg_w_42[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_3 = result_reg_w_42[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_4 = result_reg_w_42[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_5 = result_reg_w_42[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_6 = result_reg_w_42[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_7 = result_reg_w_42[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_8 = result_reg_w_42[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_9 = result_reg_w_42[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_10 = result_reg_w_42[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_11 = result_reg_w_42[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_12 = result_reg_w_42[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_13 = result_reg_w_42[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_14 = result_reg_w_42[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_15 = result_reg_w_42[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_16 = result_reg_w_42[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_17 = result_reg_w_42[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_18 = result_reg_w_42[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_19 = result_reg_w_42[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_21 = result_reg_w_42[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_22 = result_reg_w_42[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_23 = result_reg_w_42[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_24 = result_reg_w_42[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_25 = result_reg_w_42[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_26 = result_reg_w_42[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_27 = result_reg_w_42[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_28 = result_reg_w_42[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_29 = result_reg_w_42[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_30 = result_reg_w_42[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_31 = result_reg_w_42[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_32 = result_reg_w_42[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_33 = result_reg_w_42[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_34 = result_reg_w_42[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_35 = result_reg_w_42[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_36 = result_reg_w_42[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_37 = result_reg_w_42[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_38 = result_reg_w_42[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_39 = result_reg_w_42[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_40 = result_reg_w_42[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_41 = result_reg_w_42[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_42 = result_reg_w_42[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_43 = result_reg_w_42[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_44 = result_reg_w_42[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_45 = result_reg_w_42[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_46 = result_reg_w_42[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_47 = result_reg_w_42[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_48 = result_reg_w_42[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_49 = result_reg_w_42[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_50 = result_reg_w_42[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_51 = result_reg_w_42[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_52 = result_reg_w_42[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_53 = result_reg_w_42[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_54 = result_reg_w_42[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_55 = result_reg_w_42[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_56 = result_reg_w_42[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_57 = result_reg_w_42[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_58 = result_reg_w_42[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_59 = result_reg_w_42[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_60 = result_reg_w_42[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_61 = result_reg_w_42[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_62 = result_reg_w_42[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_63 = result_reg_w_42[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_64 = result_reg_w_42[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_65 = result_reg_w_42[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_66 = result_reg_w_42[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_67 = result_reg_w_42[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_68 = result_reg_w_42[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_69 = result_reg_w_42[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_70 = result_reg_w_42[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_71 = result_reg_w_42[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_72 = result_reg_w_42[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_73 = result_reg_w_42[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_74 = result_reg_w_42[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_75 = result_reg_w_42[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_76 = result_reg_w_42[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_77 = result_reg_w_42[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_78 = result_reg_w_42[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_79 = result_reg_w_42[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_80 = result_reg_w_42[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_81 = result_reg_w_42[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_82 = result_reg_w_42[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_83 = result_reg_w_42[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_84 = result_reg_w_42[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_85 = result_reg_w_42[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_86 = result_reg_w_42[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_87 = result_reg_w_42[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_88 = result_reg_w_42[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_89 = result_reg_w_42[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_90 = result_reg_w_42[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_91 = result_reg_w_42[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_92 = result_reg_w_42[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_93 = result_reg_w_42[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_94 = result_reg_w_42[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_95 = result_reg_w_42[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_96 = result_reg_w_42[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_97 = result_reg_w_42[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_98 = result_reg_w_42[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_99 = result_reg_w_42[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_100 = result_reg_w_42[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_101 = result_reg_w_42[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_102 = result_reg_w_42[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_103 = result_reg_w_42[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_104 = result_reg_w_42[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_84_105 = result_reg_w_42[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_0 = result_reg_r_42[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_1 = result_reg_r_42[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_2 = result_reg_r_42[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_3 = result_reg_r_42[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_4 = result_reg_r_42[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_5 = result_reg_r_42[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_6 = result_reg_r_42[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_7 = result_reg_r_42[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_8 = result_reg_r_42[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_9 = result_reg_r_42[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_10 = result_reg_r_42[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_11 = result_reg_r_42[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_12 = result_reg_r_42[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_13 = result_reg_r_42[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_14 = result_reg_r_42[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_15 = result_reg_r_42[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_16 = result_reg_r_42[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_17 = result_reg_r_42[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_18 = result_reg_r_42[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_20 = result_reg_r_42[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_21 = result_reg_r_42[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_22 = result_reg_r_42[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_23 = result_reg_r_42[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_24 = result_reg_r_42[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_25 = result_reg_r_42[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_26 = result_reg_r_42[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_27 = result_reg_r_42[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_28 = result_reg_r_42[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_29 = result_reg_r_42[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_30 = result_reg_r_42[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_31 = result_reg_r_42[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_32 = result_reg_r_42[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_33 = result_reg_r_42[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_34 = result_reg_r_42[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_35 = result_reg_r_42[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_36 = result_reg_r_42[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_37 = result_reg_r_42[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_38 = result_reg_r_42[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_39 = result_reg_r_42[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_40 = result_reg_r_42[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_41 = result_reg_r_42[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_42 = result_reg_r_42[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_43 = result_reg_r_42[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_44 = result_reg_r_42[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_45 = result_reg_r_42[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_46 = result_reg_r_42[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_47 = result_reg_r_42[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_48 = result_reg_r_42[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_49 = result_reg_r_42[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_50 = result_reg_r_42[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_51 = result_reg_r_42[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_52 = result_reg_r_42[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_53 = result_reg_r_42[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_54 = result_reg_r_42[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_55 = result_reg_r_42[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_56 = result_reg_r_42[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_57 = result_reg_r_42[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_58 = result_reg_r_42[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_59 = result_reg_r_42[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_60 = result_reg_r_42[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_61 = result_reg_r_42[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_62 = result_reg_r_42[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_63 = result_reg_r_42[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_64 = result_reg_r_42[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_65 = result_reg_r_42[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_66 = result_reg_r_42[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_67 = result_reg_r_42[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_68 = result_reg_r_42[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_69 = result_reg_r_42[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_70 = result_reg_r_42[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_71 = result_reg_r_42[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_72 = result_reg_r_42[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_73 = result_reg_r_42[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_74 = result_reg_r_42[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_75 = result_reg_r_42[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_76 = result_reg_r_42[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_77 = result_reg_r_42[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_78 = result_reg_r_42[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_79 = result_reg_r_42[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_80 = result_reg_r_42[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_81 = result_reg_r_42[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_82 = result_reg_r_42[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_83 = result_reg_r_42[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_84 = result_reg_r_42[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_85 = result_reg_r_42[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_86 = result_reg_r_42[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_87 = result_reg_r_42[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_88 = result_reg_r_42[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_89 = result_reg_r_42[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_90 = result_reg_r_42[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_91 = result_reg_r_42[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_92 = result_reg_r_42[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_93 = result_reg_r_42[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_94 = result_reg_r_42[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_95 = result_reg_r_42[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_96 = result_reg_r_42[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_97 = result_reg_r_42[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_98 = result_reg_r_42[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_99 = result_reg_r_42[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_100 = result_reg_r_42[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_101 = result_reg_r_42[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_102 = result_reg_r_42[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_103 = result_reg_r_42[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_104 = result_reg_r_42[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_85_105 = result_reg_r_42[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_43_hi_hi_hi_lo = {wire_res_85_98,wire_res_85_97,wire_res_85_96,wire_res_85_95,wire_res_85_94,
    wire_res_85_93,wire_res_85_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_43_hi_hi_lo_lo = {wire_res_85_84,wire_res_85_83,wire_res_85_82,wire_res_85_81,wire_res_85_80,
    wire_res_85_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_43_hi_hi_lo = {wire_res_85_91,wire_res_85_90,wire_res_85_89,wire_res_85_88,wire_res_85_87,
    wire_res_85_86,wire_res_85_85,result_reg_w_43_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_43_hi_lo_hi_lo = {wire_res_85_71,wire_res_85_70,wire_res_85_69,wire_res_85_68,wire_res_85_67,
    wire_res_85_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_43_hi_lo_lo_lo = {wire_res_85_58,wire_res_85_57,wire_res_85_56,wire_res_85_55,wire_res_85_54,
    wire_res_85_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_43_hi_lo_lo = {wire_res_85_65,wire_res_85_64,wire_res_85_63,wire_res_85_62,wire_res_85_61,
    wire_res_85_60,wire_res_85_59,result_reg_w_43_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_43_hi_lo = {wire_res_85_78,wire_res_85_77,wire_res_85_76,wire_res_85_75,wire_res_85_74,
    wire_res_85_73,wire_res_85_72,result_reg_w_43_hi_lo_hi_lo,result_reg_w_43_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_43_hi = {wire_res_85_105,wire_res_85_104,wire_res_85_103,wire_res_85_102,wire_res_85_101,
    wire_res_85_100,wire_res_85_99,result_reg_w_43_hi_hi_hi_lo,result_reg_w_43_hi_hi_lo,result_reg_w_43_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_43_lo_hi_hi_lo = {wire_res_85_45,wire_res_85_44,wire_res_85_43,wire_res_85_42,wire_res_85_41,
    wire_res_85_40,wire_res_85_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_43_lo_hi_lo_lo = {wire_res_85_31,wire_res_85_30,wire_res_85_29,wire_res_85_28,wire_res_85_27,
    wire_res_85_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_43_lo_hi_lo = {wire_res_85_38,wire_res_85_37,wire_res_85_36,wire_res_85_35,wire_res_85_34,
    wire_res_85_33,wire_res_85_32,result_reg_w_43_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [124:0] _T_11408 = {b_aux_reg_r_42, 19'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [124:0] _GEN_1314 = {{19'd0}, a_aux_reg_r_42}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_85_19 = _GEN_1314 >= _T_11408; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_43_lo_lo_hi_lo = {wire_res_85_18,wire_res_85_17,wire_res_85_16,wire_res_85_15,wire_res_85_14,
    wire_res_85_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_43_lo_lo_lo_lo = {wire_res_85_5,wire_res_85_4,wire_res_85_3,wire_res_85_2,wire_res_85_1,
    wire_res_85_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_43_lo_lo_lo = {wire_res_85_12,wire_res_85_11,wire_res_85_10,wire_res_85_9,wire_res_85_8,
    wire_res_85_7,wire_res_85_6,result_reg_w_43_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_43_lo_lo = {wire_res_85_25,wire_res_85_24,wire_res_85_23,wire_res_85_22,wire_res_85_21,
    wire_res_85_20,wire_res_85_19,result_reg_w_43_lo_lo_hi_lo,result_reg_w_43_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_43_lo = {wire_res_85_52,wire_res_85_51,wire_res_85_50,wire_res_85_49,wire_res_85_48,
    wire_res_85_47,wire_res_85_46,result_reg_w_43_lo_hi_hi_lo,result_reg_w_43_lo_hi_lo,result_reg_w_43_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_43 = {result_reg_w_43_hi,result_reg_w_43_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_86_0 = result_reg_w_43[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_1 = result_reg_w_43[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_2 = result_reg_w_43[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_3 = result_reg_w_43[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_4 = result_reg_w_43[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_5 = result_reg_w_43[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_6 = result_reg_w_43[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_7 = result_reg_w_43[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_8 = result_reg_w_43[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_9 = result_reg_w_43[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_10 = result_reg_w_43[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_11 = result_reg_w_43[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_12 = result_reg_w_43[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_13 = result_reg_w_43[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_14 = result_reg_w_43[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_15 = result_reg_w_43[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_16 = result_reg_w_43[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_17 = result_reg_w_43[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_19 = result_reg_w_43[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_20 = result_reg_w_43[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_21 = result_reg_w_43[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_22 = result_reg_w_43[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_23 = result_reg_w_43[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_24 = result_reg_w_43[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_25 = result_reg_w_43[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_26 = result_reg_w_43[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_27 = result_reg_w_43[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_28 = result_reg_w_43[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_29 = result_reg_w_43[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_30 = result_reg_w_43[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_31 = result_reg_w_43[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_32 = result_reg_w_43[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_33 = result_reg_w_43[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_34 = result_reg_w_43[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_35 = result_reg_w_43[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_36 = result_reg_w_43[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_37 = result_reg_w_43[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_38 = result_reg_w_43[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_39 = result_reg_w_43[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_40 = result_reg_w_43[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_41 = result_reg_w_43[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_42 = result_reg_w_43[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_43 = result_reg_w_43[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_44 = result_reg_w_43[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_45 = result_reg_w_43[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_46 = result_reg_w_43[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_47 = result_reg_w_43[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_48 = result_reg_w_43[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_49 = result_reg_w_43[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_50 = result_reg_w_43[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_51 = result_reg_w_43[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_52 = result_reg_w_43[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_53 = result_reg_w_43[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_54 = result_reg_w_43[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_55 = result_reg_w_43[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_56 = result_reg_w_43[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_57 = result_reg_w_43[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_58 = result_reg_w_43[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_59 = result_reg_w_43[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_60 = result_reg_w_43[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_61 = result_reg_w_43[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_62 = result_reg_w_43[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_63 = result_reg_w_43[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_64 = result_reg_w_43[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_65 = result_reg_w_43[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_66 = result_reg_w_43[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_67 = result_reg_w_43[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_68 = result_reg_w_43[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_69 = result_reg_w_43[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_70 = result_reg_w_43[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_71 = result_reg_w_43[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_72 = result_reg_w_43[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_73 = result_reg_w_43[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_74 = result_reg_w_43[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_75 = result_reg_w_43[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_76 = result_reg_w_43[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_77 = result_reg_w_43[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_78 = result_reg_w_43[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_79 = result_reg_w_43[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_80 = result_reg_w_43[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_81 = result_reg_w_43[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_82 = result_reg_w_43[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_83 = result_reg_w_43[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_84 = result_reg_w_43[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_85 = result_reg_w_43[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_86 = result_reg_w_43[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_87 = result_reg_w_43[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_88 = result_reg_w_43[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_89 = result_reg_w_43[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_90 = result_reg_w_43[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_91 = result_reg_w_43[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_92 = result_reg_w_43[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_93 = result_reg_w_43[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_94 = result_reg_w_43[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_95 = result_reg_w_43[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_96 = result_reg_w_43[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_97 = result_reg_w_43[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_98 = result_reg_w_43[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_99 = result_reg_w_43[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_100 = result_reg_w_43[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_101 = result_reg_w_43[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_102 = result_reg_w_43[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_103 = result_reg_w_43[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_104 = result_reg_w_43[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_86_105 = result_reg_w_43[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_0 = result_reg_r_43[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_1 = result_reg_r_43[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_2 = result_reg_r_43[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_3 = result_reg_r_43[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_4 = result_reg_r_43[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_5 = result_reg_r_43[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_6 = result_reg_r_43[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_7 = result_reg_r_43[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_8 = result_reg_r_43[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_9 = result_reg_r_43[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_10 = result_reg_r_43[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_11 = result_reg_r_43[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_12 = result_reg_r_43[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_13 = result_reg_r_43[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_14 = result_reg_r_43[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_15 = result_reg_r_43[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_16 = result_reg_r_43[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_18 = result_reg_r_43[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_19 = result_reg_r_43[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_20 = result_reg_r_43[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_21 = result_reg_r_43[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_22 = result_reg_r_43[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_23 = result_reg_r_43[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_24 = result_reg_r_43[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_25 = result_reg_r_43[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_26 = result_reg_r_43[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_27 = result_reg_r_43[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_28 = result_reg_r_43[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_29 = result_reg_r_43[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_30 = result_reg_r_43[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_31 = result_reg_r_43[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_32 = result_reg_r_43[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_33 = result_reg_r_43[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_34 = result_reg_r_43[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_35 = result_reg_r_43[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_36 = result_reg_r_43[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_37 = result_reg_r_43[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_38 = result_reg_r_43[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_39 = result_reg_r_43[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_40 = result_reg_r_43[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_41 = result_reg_r_43[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_42 = result_reg_r_43[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_43 = result_reg_r_43[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_44 = result_reg_r_43[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_45 = result_reg_r_43[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_46 = result_reg_r_43[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_47 = result_reg_r_43[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_48 = result_reg_r_43[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_49 = result_reg_r_43[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_50 = result_reg_r_43[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_51 = result_reg_r_43[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_52 = result_reg_r_43[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_53 = result_reg_r_43[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_54 = result_reg_r_43[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_55 = result_reg_r_43[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_56 = result_reg_r_43[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_57 = result_reg_r_43[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_58 = result_reg_r_43[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_59 = result_reg_r_43[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_60 = result_reg_r_43[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_61 = result_reg_r_43[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_62 = result_reg_r_43[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_63 = result_reg_r_43[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_64 = result_reg_r_43[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_65 = result_reg_r_43[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_66 = result_reg_r_43[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_67 = result_reg_r_43[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_68 = result_reg_r_43[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_69 = result_reg_r_43[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_70 = result_reg_r_43[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_71 = result_reg_r_43[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_72 = result_reg_r_43[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_73 = result_reg_r_43[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_74 = result_reg_r_43[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_75 = result_reg_r_43[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_76 = result_reg_r_43[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_77 = result_reg_r_43[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_78 = result_reg_r_43[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_79 = result_reg_r_43[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_80 = result_reg_r_43[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_81 = result_reg_r_43[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_82 = result_reg_r_43[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_83 = result_reg_r_43[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_84 = result_reg_r_43[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_85 = result_reg_r_43[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_86 = result_reg_r_43[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_87 = result_reg_r_43[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_88 = result_reg_r_43[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_89 = result_reg_r_43[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_90 = result_reg_r_43[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_91 = result_reg_r_43[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_92 = result_reg_r_43[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_93 = result_reg_r_43[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_94 = result_reg_r_43[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_95 = result_reg_r_43[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_96 = result_reg_r_43[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_97 = result_reg_r_43[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_98 = result_reg_r_43[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_99 = result_reg_r_43[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_100 = result_reg_r_43[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_101 = result_reg_r_43[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_102 = result_reg_r_43[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_103 = result_reg_r_43[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_104 = result_reg_r_43[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_87_105 = result_reg_r_43[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_44_hi_hi_hi_lo = {wire_res_87_98,wire_res_87_97,wire_res_87_96,wire_res_87_95,wire_res_87_94,
    wire_res_87_93,wire_res_87_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_44_hi_hi_lo_lo = {wire_res_87_84,wire_res_87_83,wire_res_87_82,wire_res_87_81,wire_res_87_80,
    wire_res_87_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_44_hi_hi_lo = {wire_res_87_91,wire_res_87_90,wire_res_87_89,wire_res_87_88,wire_res_87_87,
    wire_res_87_86,wire_res_87_85,result_reg_w_44_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_44_hi_lo_hi_lo = {wire_res_87_71,wire_res_87_70,wire_res_87_69,wire_res_87_68,wire_res_87_67,
    wire_res_87_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_44_hi_lo_lo_lo = {wire_res_87_58,wire_res_87_57,wire_res_87_56,wire_res_87_55,wire_res_87_54,
    wire_res_87_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_44_hi_lo_lo = {wire_res_87_65,wire_res_87_64,wire_res_87_63,wire_res_87_62,wire_res_87_61,
    wire_res_87_60,wire_res_87_59,result_reg_w_44_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_44_hi_lo = {wire_res_87_78,wire_res_87_77,wire_res_87_76,wire_res_87_75,wire_res_87_74,
    wire_res_87_73,wire_res_87_72,result_reg_w_44_hi_lo_hi_lo,result_reg_w_44_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_44_hi = {wire_res_87_105,wire_res_87_104,wire_res_87_103,wire_res_87_102,wire_res_87_101,
    wire_res_87_100,wire_res_87_99,result_reg_w_44_hi_hi_hi_lo,result_reg_w_44_hi_hi_lo,result_reg_w_44_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_44_lo_hi_hi_lo = {wire_res_87_45,wire_res_87_44,wire_res_87_43,wire_res_87_42,wire_res_87_41,
    wire_res_87_40,wire_res_87_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_44_lo_hi_lo_lo = {wire_res_87_31,wire_res_87_30,wire_res_87_29,wire_res_87_28,wire_res_87_27,
    wire_res_87_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_44_lo_hi_lo = {wire_res_87_38,wire_res_87_37,wire_res_87_36,wire_res_87_35,wire_res_87_34,
    wire_res_87_33,wire_res_87_32,result_reg_w_44_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [122:0] _T_11412 = {b_aux_reg_r_43, 17'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [122:0] _GEN_1315 = {{17'd0}, a_aux_reg_r_43}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_87_17 = _GEN_1315 >= _T_11412; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_44_lo_lo_hi_lo = {wire_res_87_18,wire_res_87_17,wire_res_87_16,wire_res_87_15,wire_res_87_14,
    wire_res_87_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_44_lo_lo_lo_lo = {wire_res_87_5,wire_res_87_4,wire_res_87_3,wire_res_87_2,wire_res_87_1,
    wire_res_87_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_44_lo_lo_lo = {wire_res_87_12,wire_res_87_11,wire_res_87_10,wire_res_87_9,wire_res_87_8,
    wire_res_87_7,wire_res_87_6,result_reg_w_44_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_44_lo_lo = {wire_res_87_25,wire_res_87_24,wire_res_87_23,wire_res_87_22,wire_res_87_21,
    wire_res_87_20,wire_res_87_19,result_reg_w_44_lo_lo_hi_lo,result_reg_w_44_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_44_lo = {wire_res_87_52,wire_res_87_51,wire_res_87_50,wire_res_87_49,wire_res_87_48,
    wire_res_87_47,wire_res_87_46,result_reg_w_44_lo_hi_hi_lo,result_reg_w_44_lo_hi_lo,result_reg_w_44_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_44 = {result_reg_w_44_hi,result_reg_w_44_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_88_0 = result_reg_w_44[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_1 = result_reg_w_44[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_2 = result_reg_w_44[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_3 = result_reg_w_44[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_4 = result_reg_w_44[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_5 = result_reg_w_44[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_6 = result_reg_w_44[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_7 = result_reg_w_44[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_8 = result_reg_w_44[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_9 = result_reg_w_44[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_10 = result_reg_w_44[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_11 = result_reg_w_44[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_12 = result_reg_w_44[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_13 = result_reg_w_44[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_14 = result_reg_w_44[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_15 = result_reg_w_44[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_17 = result_reg_w_44[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_18 = result_reg_w_44[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_19 = result_reg_w_44[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_20 = result_reg_w_44[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_21 = result_reg_w_44[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_22 = result_reg_w_44[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_23 = result_reg_w_44[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_24 = result_reg_w_44[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_25 = result_reg_w_44[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_26 = result_reg_w_44[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_27 = result_reg_w_44[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_28 = result_reg_w_44[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_29 = result_reg_w_44[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_30 = result_reg_w_44[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_31 = result_reg_w_44[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_32 = result_reg_w_44[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_33 = result_reg_w_44[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_34 = result_reg_w_44[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_35 = result_reg_w_44[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_36 = result_reg_w_44[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_37 = result_reg_w_44[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_38 = result_reg_w_44[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_39 = result_reg_w_44[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_40 = result_reg_w_44[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_41 = result_reg_w_44[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_42 = result_reg_w_44[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_43 = result_reg_w_44[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_44 = result_reg_w_44[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_45 = result_reg_w_44[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_46 = result_reg_w_44[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_47 = result_reg_w_44[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_48 = result_reg_w_44[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_49 = result_reg_w_44[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_50 = result_reg_w_44[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_51 = result_reg_w_44[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_52 = result_reg_w_44[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_53 = result_reg_w_44[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_54 = result_reg_w_44[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_55 = result_reg_w_44[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_56 = result_reg_w_44[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_57 = result_reg_w_44[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_58 = result_reg_w_44[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_59 = result_reg_w_44[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_60 = result_reg_w_44[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_61 = result_reg_w_44[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_62 = result_reg_w_44[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_63 = result_reg_w_44[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_64 = result_reg_w_44[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_65 = result_reg_w_44[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_66 = result_reg_w_44[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_67 = result_reg_w_44[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_68 = result_reg_w_44[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_69 = result_reg_w_44[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_70 = result_reg_w_44[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_71 = result_reg_w_44[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_72 = result_reg_w_44[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_73 = result_reg_w_44[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_74 = result_reg_w_44[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_75 = result_reg_w_44[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_76 = result_reg_w_44[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_77 = result_reg_w_44[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_78 = result_reg_w_44[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_79 = result_reg_w_44[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_80 = result_reg_w_44[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_81 = result_reg_w_44[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_82 = result_reg_w_44[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_83 = result_reg_w_44[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_84 = result_reg_w_44[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_85 = result_reg_w_44[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_86 = result_reg_w_44[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_87 = result_reg_w_44[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_88 = result_reg_w_44[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_89 = result_reg_w_44[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_90 = result_reg_w_44[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_91 = result_reg_w_44[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_92 = result_reg_w_44[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_93 = result_reg_w_44[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_94 = result_reg_w_44[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_95 = result_reg_w_44[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_96 = result_reg_w_44[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_97 = result_reg_w_44[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_98 = result_reg_w_44[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_99 = result_reg_w_44[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_100 = result_reg_w_44[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_101 = result_reg_w_44[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_102 = result_reg_w_44[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_103 = result_reg_w_44[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_104 = result_reg_w_44[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_88_105 = result_reg_w_44[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_0 = result_reg_r_44[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_1 = result_reg_r_44[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_2 = result_reg_r_44[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_3 = result_reg_r_44[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_4 = result_reg_r_44[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_5 = result_reg_r_44[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_6 = result_reg_r_44[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_7 = result_reg_r_44[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_8 = result_reg_r_44[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_9 = result_reg_r_44[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_10 = result_reg_r_44[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_11 = result_reg_r_44[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_12 = result_reg_r_44[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_13 = result_reg_r_44[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_14 = result_reg_r_44[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_16 = result_reg_r_44[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_17 = result_reg_r_44[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_18 = result_reg_r_44[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_19 = result_reg_r_44[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_20 = result_reg_r_44[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_21 = result_reg_r_44[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_22 = result_reg_r_44[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_23 = result_reg_r_44[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_24 = result_reg_r_44[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_25 = result_reg_r_44[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_26 = result_reg_r_44[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_27 = result_reg_r_44[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_28 = result_reg_r_44[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_29 = result_reg_r_44[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_30 = result_reg_r_44[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_31 = result_reg_r_44[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_32 = result_reg_r_44[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_33 = result_reg_r_44[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_34 = result_reg_r_44[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_35 = result_reg_r_44[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_36 = result_reg_r_44[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_37 = result_reg_r_44[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_38 = result_reg_r_44[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_39 = result_reg_r_44[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_40 = result_reg_r_44[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_41 = result_reg_r_44[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_42 = result_reg_r_44[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_43 = result_reg_r_44[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_44 = result_reg_r_44[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_45 = result_reg_r_44[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_46 = result_reg_r_44[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_47 = result_reg_r_44[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_48 = result_reg_r_44[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_49 = result_reg_r_44[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_50 = result_reg_r_44[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_51 = result_reg_r_44[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_52 = result_reg_r_44[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_53 = result_reg_r_44[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_54 = result_reg_r_44[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_55 = result_reg_r_44[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_56 = result_reg_r_44[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_57 = result_reg_r_44[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_58 = result_reg_r_44[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_59 = result_reg_r_44[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_60 = result_reg_r_44[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_61 = result_reg_r_44[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_62 = result_reg_r_44[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_63 = result_reg_r_44[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_64 = result_reg_r_44[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_65 = result_reg_r_44[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_66 = result_reg_r_44[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_67 = result_reg_r_44[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_68 = result_reg_r_44[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_69 = result_reg_r_44[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_70 = result_reg_r_44[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_71 = result_reg_r_44[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_72 = result_reg_r_44[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_73 = result_reg_r_44[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_74 = result_reg_r_44[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_75 = result_reg_r_44[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_76 = result_reg_r_44[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_77 = result_reg_r_44[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_78 = result_reg_r_44[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_79 = result_reg_r_44[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_80 = result_reg_r_44[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_81 = result_reg_r_44[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_82 = result_reg_r_44[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_83 = result_reg_r_44[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_84 = result_reg_r_44[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_85 = result_reg_r_44[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_86 = result_reg_r_44[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_87 = result_reg_r_44[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_88 = result_reg_r_44[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_89 = result_reg_r_44[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_90 = result_reg_r_44[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_91 = result_reg_r_44[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_92 = result_reg_r_44[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_93 = result_reg_r_44[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_94 = result_reg_r_44[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_95 = result_reg_r_44[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_96 = result_reg_r_44[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_97 = result_reg_r_44[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_98 = result_reg_r_44[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_99 = result_reg_r_44[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_100 = result_reg_r_44[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_101 = result_reg_r_44[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_102 = result_reg_r_44[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_103 = result_reg_r_44[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_104 = result_reg_r_44[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_89_105 = result_reg_r_44[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_45_hi_hi_hi_lo = {wire_res_89_98,wire_res_89_97,wire_res_89_96,wire_res_89_95,wire_res_89_94,
    wire_res_89_93,wire_res_89_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_45_hi_hi_lo_lo = {wire_res_89_84,wire_res_89_83,wire_res_89_82,wire_res_89_81,wire_res_89_80,
    wire_res_89_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_45_hi_hi_lo = {wire_res_89_91,wire_res_89_90,wire_res_89_89,wire_res_89_88,wire_res_89_87,
    wire_res_89_86,wire_res_89_85,result_reg_w_45_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_45_hi_lo_hi_lo = {wire_res_89_71,wire_res_89_70,wire_res_89_69,wire_res_89_68,wire_res_89_67,
    wire_res_89_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_45_hi_lo_lo_lo = {wire_res_89_58,wire_res_89_57,wire_res_89_56,wire_res_89_55,wire_res_89_54,
    wire_res_89_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_45_hi_lo_lo = {wire_res_89_65,wire_res_89_64,wire_res_89_63,wire_res_89_62,wire_res_89_61,
    wire_res_89_60,wire_res_89_59,result_reg_w_45_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_45_hi_lo = {wire_res_89_78,wire_res_89_77,wire_res_89_76,wire_res_89_75,wire_res_89_74,
    wire_res_89_73,wire_res_89_72,result_reg_w_45_hi_lo_hi_lo,result_reg_w_45_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_45_hi = {wire_res_89_105,wire_res_89_104,wire_res_89_103,wire_res_89_102,wire_res_89_101,
    wire_res_89_100,wire_res_89_99,result_reg_w_45_hi_hi_hi_lo,result_reg_w_45_hi_hi_lo,result_reg_w_45_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_45_lo_hi_hi_lo = {wire_res_89_45,wire_res_89_44,wire_res_89_43,wire_res_89_42,wire_res_89_41,
    wire_res_89_40,wire_res_89_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_45_lo_hi_lo_lo = {wire_res_89_31,wire_res_89_30,wire_res_89_29,wire_res_89_28,wire_res_89_27,
    wire_res_89_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_45_lo_hi_lo = {wire_res_89_38,wire_res_89_37,wire_res_89_36,wire_res_89_35,wire_res_89_34,
    wire_res_89_33,wire_res_89_32,result_reg_w_45_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [120:0] _T_11416 = {b_aux_reg_r_44, 15'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [120:0] _GEN_1316 = {{15'd0}, a_aux_reg_r_44}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_89_15 = _GEN_1316 >= _T_11416; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_45_lo_lo_hi_lo = {wire_res_89_18,wire_res_89_17,wire_res_89_16,wire_res_89_15,wire_res_89_14,
    wire_res_89_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_45_lo_lo_lo_lo = {wire_res_89_5,wire_res_89_4,wire_res_89_3,wire_res_89_2,wire_res_89_1,
    wire_res_89_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_45_lo_lo_lo = {wire_res_89_12,wire_res_89_11,wire_res_89_10,wire_res_89_9,wire_res_89_8,
    wire_res_89_7,wire_res_89_6,result_reg_w_45_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_45_lo_lo = {wire_res_89_25,wire_res_89_24,wire_res_89_23,wire_res_89_22,wire_res_89_21,
    wire_res_89_20,wire_res_89_19,result_reg_w_45_lo_lo_hi_lo,result_reg_w_45_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_45_lo = {wire_res_89_52,wire_res_89_51,wire_res_89_50,wire_res_89_49,wire_res_89_48,
    wire_res_89_47,wire_res_89_46,result_reg_w_45_lo_hi_hi_lo,result_reg_w_45_lo_hi_lo,result_reg_w_45_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_45 = {result_reg_w_45_hi,result_reg_w_45_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_90_0 = result_reg_w_45[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_1 = result_reg_w_45[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_2 = result_reg_w_45[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_3 = result_reg_w_45[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_4 = result_reg_w_45[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_5 = result_reg_w_45[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_6 = result_reg_w_45[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_7 = result_reg_w_45[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_8 = result_reg_w_45[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_9 = result_reg_w_45[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_10 = result_reg_w_45[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_11 = result_reg_w_45[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_12 = result_reg_w_45[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_13 = result_reg_w_45[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_15 = result_reg_w_45[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_16 = result_reg_w_45[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_17 = result_reg_w_45[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_18 = result_reg_w_45[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_19 = result_reg_w_45[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_20 = result_reg_w_45[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_21 = result_reg_w_45[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_22 = result_reg_w_45[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_23 = result_reg_w_45[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_24 = result_reg_w_45[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_25 = result_reg_w_45[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_26 = result_reg_w_45[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_27 = result_reg_w_45[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_28 = result_reg_w_45[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_29 = result_reg_w_45[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_30 = result_reg_w_45[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_31 = result_reg_w_45[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_32 = result_reg_w_45[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_33 = result_reg_w_45[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_34 = result_reg_w_45[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_35 = result_reg_w_45[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_36 = result_reg_w_45[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_37 = result_reg_w_45[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_38 = result_reg_w_45[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_39 = result_reg_w_45[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_40 = result_reg_w_45[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_41 = result_reg_w_45[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_42 = result_reg_w_45[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_43 = result_reg_w_45[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_44 = result_reg_w_45[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_45 = result_reg_w_45[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_46 = result_reg_w_45[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_47 = result_reg_w_45[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_48 = result_reg_w_45[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_49 = result_reg_w_45[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_50 = result_reg_w_45[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_51 = result_reg_w_45[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_52 = result_reg_w_45[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_53 = result_reg_w_45[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_54 = result_reg_w_45[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_55 = result_reg_w_45[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_56 = result_reg_w_45[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_57 = result_reg_w_45[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_58 = result_reg_w_45[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_59 = result_reg_w_45[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_60 = result_reg_w_45[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_61 = result_reg_w_45[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_62 = result_reg_w_45[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_63 = result_reg_w_45[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_64 = result_reg_w_45[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_65 = result_reg_w_45[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_66 = result_reg_w_45[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_67 = result_reg_w_45[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_68 = result_reg_w_45[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_69 = result_reg_w_45[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_70 = result_reg_w_45[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_71 = result_reg_w_45[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_72 = result_reg_w_45[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_73 = result_reg_w_45[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_74 = result_reg_w_45[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_75 = result_reg_w_45[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_76 = result_reg_w_45[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_77 = result_reg_w_45[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_78 = result_reg_w_45[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_79 = result_reg_w_45[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_80 = result_reg_w_45[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_81 = result_reg_w_45[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_82 = result_reg_w_45[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_83 = result_reg_w_45[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_84 = result_reg_w_45[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_85 = result_reg_w_45[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_86 = result_reg_w_45[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_87 = result_reg_w_45[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_88 = result_reg_w_45[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_89 = result_reg_w_45[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_90 = result_reg_w_45[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_91 = result_reg_w_45[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_92 = result_reg_w_45[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_93 = result_reg_w_45[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_94 = result_reg_w_45[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_95 = result_reg_w_45[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_96 = result_reg_w_45[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_97 = result_reg_w_45[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_98 = result_reg_w_45[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_99 = result_reg_w_45[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_100 = result_reg_w_45[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_101 = result_reg_w_45[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_102 = result_reg_w_45[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_103 = result_reg_w_45[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_104 = result_reg_w_45[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_90_105 = result_reg_w_45[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_0 = result_reg_r_45[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_1 = result_reg_r_45[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_2 = result_reg_r_45[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_3 = result_reg_r_45[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_4 = result_reg_r_45[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_5 = result_reg_r_45[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_6 = result_reg_r_45[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_7 = result_reg_r_45[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_8 = result_reg_r_45[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_9 = result_reg_r_45[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_10 = result_reg_r_45[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_11 = result_reg_r_45[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_12 = result_reg_r_45[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_14 = result_reg_r_45[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_15 = result_reg_r_45[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_16 = result_reg_r_45[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_17 = result_reg_r_45[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_18 = result_reg_r_45[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_19 = result_reg_r_45[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_20 = result_reg_r_45[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_21 = result_reg_r_45[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_22 = result_reg_r_45[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_23 = result_reg_r_45[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_24 = result_reg_r_45[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_25 = result_reg_r_45[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_26 = result_reg_r_45[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_27 = result_reg_r_45[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_28 = result_reg_r_45[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_29 = result_reg_r_45[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_30 = result_reg_r_45[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_31 = result_reg_r_45[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_32 = result_reg_r_45[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_33 = result_reg_r_45[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_34 = result_reg_r_45[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_35 = result_reg_r_45[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_36 = result_reg_r_45[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_37 = result_reg_r_45[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_38 = result_reg_r_45[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_39 = result_reg_r_45[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_40 = result_reg_r_45[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_41 = result_reg_r_45[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_42 = result_reg_r_45[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_43 = result_reg_r_45[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_44 = result_reg_r_45[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_45 = result_reg_r_45[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_46 = result_reg_r_45[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_47 = result_reg_r_45[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_48 = result_reg_r_45[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_49 = result_reg_r_45[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_50 = result_reg_r_45[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_51 = result_reg_r_45[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_52 = result_reg_r_45[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_53 = result_reg_r_45[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_54 = result_reg_r_45[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_55 = result_reg_r_45[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_56 = result_reg_r_45[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_57 = result_reg_r_45[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_58 = result_reg_r_45[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_59 = result_reg_r_45[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_60 = result_reg_r_45[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_61 = result_reg_r_45[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_62 = result_reg_r_45[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_63 = result_reg_r_45[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_64 = result_reg_r_45[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_65 = result_reg_r_45[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_66 = result_reg_r_45[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_67 = result_reg_r_45[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_68 = result_reg_r_45[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_69 = result_reg_r_45[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_70 = result_reg_r_45[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_71 = result_reg_r_45[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_72 = result_reg_r_45[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_73 = result_reg_r_45[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_74 = result_reg_r_45[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_75 = result_reg_r_45[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_76 = result_reg_r_45[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_77 = result_reg_r_45[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_78 = result_reg_r_45[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_79 = result_reg_r_45[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_80 = result_reg_r_45[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_81 = result_reg_r_45[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_82 = result_reg_r_45[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_83 = result_reg_r_45[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_84 = result_reg_r_45[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_85 = result_reg_r_45[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_86 = result_reg_r_45[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_87 = result_reg_r_45[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_88 = result_reg_r_45[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_89 = result_reg_r_45[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_90 = result_reg_r_45[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_91 = result_reg_r_45[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_92 = result_reg_r_45[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_93 = result_reg_r_45[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_94 = result_reg_r_45[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_95 = result_reg_r_45[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_96 = result_reg_r_45[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_97 = result_reg_r_45[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_98 = result_reg_r_45[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_99 = result_reg_r_45[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_100 = result_reg_r_45[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_101 = result_reg_r_45[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_102 = result_reg_r_45[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_103 = result_reg_r_45[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_104 = result_reg_r_45[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_91_105 = result_reg_r_45[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_46_hi_hi_hi_lo = {wire_res_91_98,wire_res_91_97,wire_res_91_96,wire_res_91_95,wire_res_91_94,
    wire_res_91_93,wire_res_91_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_46_hi_hi_lo_lo = {wire_res_91_84,wire_res_91_83,wire_res_91_82,wire_res_91_81,wire_res_91_80,
    wire_res_91_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_46_hi_hi_lo = {wire_res_91_91,wire_res_91_90,wire_res_91_89,wire_res_91_88,wire_res_91_87,
    wire_res_91_86,wire_res_91_85,result_reg_w_46_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_46_hi_lo_hi_lo = {wire_res_91_71,wire_res_91_70,wire_res_91_69,wire_res_91_68,wire_res_91_67,
    wire_res_91_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_46_hi_lo_lo_lo = {wire_res_91_58,wire_res_91_57,wire_res_91_56,wire_res_91_55,wire_res_91_54,
    wire_res_91_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_46_hi_lo_lo = {wire_res_91_65,wire_res_91_64,wire_res_91_63,wire_res_91_62,wire_res_91_61,
    wire_res_91_60,wire_res_91_59,result_reg_w_46_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_46_hi_lo = {wire_res_91_78,wire_res_91_77,wire_res_91_76,wire_res_91_75,wire_res_91_74,
    wire_res_91_73,wire_res_91_72,result_reg_w_46_hi_lo_hi_lo,result_reg_w_46_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_46_hi = {wire_res_91_105,wire_res_91_104,wire_res_91_103,wire_res_91_102,wire_res_91_101,
    wire_res_91_100,wire_res_91_99,result_reg_w_46_hi_hi_hi_lo,result_reg_w_46_hi_hi_lo,result_reg_w_46_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_46_lo_hi_hi_lo = {wire_res_91_45,wire_res_91_44,wire_res_91_43,wire_res_91_42,wire_res_91_41,
    wire_res_91_40,wire_res_91_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_46_lo_hi_lo_lo = {wire_res_91_31,wire_res_91_30,wire_res_91_29,wire_res_91_28,wire_res_91_27,
    wire_res_91_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_46_lo_hi_lo = {wire_res_91_38,wire_res_91_37,wire_res_91_36,wire_res_91_35,wire_res_91_34,
    wire_res_91_33,wire_res_91_32,result_reg_w_46_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [118:0] _T_11420 = {b_aux_reg_r_45, 13'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [118:0] _GEN_1317 = {{13'd0}, a_aux_reg_r_45}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_91_13 = _GEN_1317 >= _T_11420; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_46_lo_lo_hi_lo = {wire_res_91_18,wire_res_91_17,wire_res_91_16,wire_res_91_15,wire_res_91_14,
    wire_res_91_13}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_46_lo_lo_lo_lo = {wire_res_91_5,wire_res_91_4,wire_res_91_3,wire_res_91_2,wire_res_91_1,
    wire_res_91_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_46_lo_lo_lo = {wire_res_91_12,wire_res_91_11,wire_res_91_10,wire_res_91_9,wire_res_91_8,
    wire_res_91_7,wire_res_91_6,result_reg_w_46_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_46_lo_lo = {wire_res_91_25,wire_res_91_24,wire_res_91_23,wire_res_91_22,wire_res_91_21,
    wire_res_91_20,wire_res_91_19,result_reg_w_46_lo_lo_hi_lo,result_reg_w_46_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_46_lo = {wire_res_91_52,wire_res_91_51,wire_res_91_50,wire_res_91_49,wire_res_91_48,
    wire_res_91_47,wire_res_91_46,result_reg_w_46_lo_hi_hi_lo,result_reg_w_46_lo_hi_lo,result_reg_w_46_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_46 = {result_reg_w_46_hi,result_reg_w_46_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_92_0 = result_reg_w_46[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_1 = result_reg_w_46[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_2 = result_reg_w_46[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_3 = result_reg_w_46[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_4 = result_reg_w_46[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_5 = result_reg_w_46[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_6 = result_reg_w_46[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_7 = result_reg_w_46[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_8 = result_reg_w_46[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_9 = result_reg_w_46[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_10 = result_reg_w_46[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_11 = result_reg_w_46[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_13 = result_reg_w_46[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_14 = result_reg_w_46[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_15 = result_reg_w_46[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_16 = result_reg_w_46[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_17 = result_reg_w_46[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_18 = result_reg_w_46[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_19 = result_reg_w_46[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_20 = result_reg_w_46[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_21 = result_reg_w_46[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_22 = result_reg_w_46[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_23 = result_reg_w_46[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_24 = result_reg_w_46[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_25 = result_reg_w_46[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_26 = result_reg_w_46[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_27 = result_reg_w_46[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_28 = result_reg_w_46[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_29 = result_reg_w_46[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_30 = result_reg_w_46[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_31 = result_reg_w_46[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_32 = result_reg_w_46[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_33 = result_reg_w_46[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_34 = result_reg_w_46[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_35 = result_reg_w_46[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_36 = result_reg_w_46[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_37 = result_reg_w_46[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_38 = result_reg_w_46[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_39 = result_reg_w_46[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_40 = result_reg_w_46[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_41 = result_reg_w_46[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_42 = result_reg_w_46[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_43 = result_reg_w_46[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_44 = result_reg_w_46[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_45 = result_reg_w_46[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_46 = result_reg_w_46[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_47 = result_reg_w_46[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_48 = result_reg_w_46[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_49 = result_reg_w_46[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_50 = result_reg_w_46[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_51 = result_reg_w_46[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_52 = result_reg_w_46[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_53 = result_reg_w_46[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_54 = result_reg_w_46[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_55 = result_reg_w_46[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_56 = result_reg_w_46[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_57 = result_reg_w_46[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_58 = result_reg_w_46[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_59 = result_reg_w_46[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_60 = result_reg_w_46[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_61 = result_reg_w_46[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_62 = result_reg_w_46[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_63 = result_reg_w_46[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_64 = result_reg_w_46[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_65 = result_reg_w_46[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_66 = result_reg_w_46[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_67 = result_reg_w_46[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_68 = result_reg_w_46[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_69 = result_reg_w_46[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_70 = result_reg_w_46[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_71 = result_reg_w_46[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_72 = result_reg_w_46[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_73 = result_reg_w_46[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_74 = result_reg_w_46[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_75 = result_reg_w_46[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_76 = result_reg_w_46[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_77 = result_reg_w_46[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_78 = result_reg_w_46[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_79 = result_reg_w_46[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_80 = result_reg_w_46[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_81 = result_reg_w_46[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_82 = result_reg_w_46[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_83 = result_reg_w_46[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_84 = result_reg_w_46[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_85 = result_reg_w_46[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_86 = result_reg_w_46[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_87 = result_reg_w_46[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_88 = result_reg_w_46[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_89 = result_reg_w_46[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_90 = result_reg_w_46[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_91 = result_reg_w_46[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_92 = result_reg_w_46[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_93 = result_reg_w_46[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_94 = result_reg_w_46[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_95 = result_reg_w_46[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_96 = result_reg_w_46[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_97 = result_reg_w_46[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_98 = result_reg_w_46[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_99 = result_reg_w_46[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_100 = result_reg_w_46[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_101 = result_reg_w_46[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_102 = result_reg_w_46[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_103 = result_reg_w_46[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_104 = result_reg_w_46[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_92_105 = result_reg_w_46[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_0 = result_reg_r_46[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_1 = result_reg_r_46[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_2 = result_reg_r_46[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_3 = result_reg_r_46[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_4 = result_reg_r_46[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_5 = result_reg_r_46[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_6 = result_reg_r_46[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_7 = result_reg_r_46[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_8 = result_reg_r_46[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_9 = result_reg_r_46[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_10 = result_reg_r_46[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_12 = result_reg_r_46[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_13 = result_reg_r_46[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_14 = result_reg_r_46[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_15 = result_reg_r_46[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_16 = result_reg_r_46[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_17 = result_reg_r_46[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_18 = result_reg_r_46[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_19 = result_reg_r_46[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_20 = result_reg_r_46[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_21 = result_reg_r_46[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_22 = result_reg_r_46[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_23 = result_reg_r_46[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_24 = result_reg_r_46[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_25 = result_reg_r_46[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_26 = result_reg_r_46[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_27 = result_reg_r_46[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_28 = result_reg_r_46[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_29 = result_reg_r_46[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_30 = result_reg_r_46[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_31 = result_reg_r_46[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_32 = result_reg_r_46[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_33 = result_reg_r_46[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_34 = result_reg_r_46[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_35 = result_reg_r_46[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_36 = result_reg_r_46[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_37 = result_reg_r_46[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_38 = result_reg_r_46[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_39 = result_reg_r_46[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_40 = result_reg_r_46[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_41 = result_reg_r_46[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_42 = result_reg_r_46[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_43 = result_reg_r_46[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_44 = result_reg_r_46[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_45 = result_reg_r_46[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_46 = result_reg_r_46[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_47 = result_reg_r_46[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_48 = result_reg_r_46[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_49 = result_reg_r_46[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_50 = result_reg_r_46[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_51 = result_reg_r_46[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_52 = result_reg_r_46[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_53 = result_reg_r_46[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_54 = result_reg_r_46[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_55 = result_reg_r_46[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_56 = result_reg_r_46[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_57 = result_reg_r_46[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_58 = result_reg_r_46[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_59 = result_reg_r_46[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_60 = result_reg_r_46[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_61 = result_reg_r_46[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_62 = result_reg_r_46[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_63 = result_reg_r_46[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_64 = result_reg_r_46[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_65 = result_reg_r_46[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_66 = result_reg_r_46[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_67 = result_reg_r_46[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_68 = result_reg_r_46[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_69 = result_reg_r_46[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_70 = result_reg_r_46[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_71 = result_reg_r_46[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_72 = result_reg_r_46[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_73 = result_reg_r_46[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_74 = result_reg_r_46[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_75 = result_reg_r_46[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_76 = result_reg_r_46[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_77 = result_reg_r_46[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_78 = result_reg_r_46[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_79 = result_reg_r_46[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_80 = result_reg_r_46[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_81 = result_reg_r_46[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_82 = result_reg_r_46[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_83 = result_reg_r_46[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_84 = result_reg_r_46[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_85 = result_reg_r_46[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_86 = result_reg_r_46[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_87 = result_reg_r_46[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_88 = result_reg_r_46[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_89 = result_reg_r_46[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_90 = result_reg_r_46[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_91 = result_reg_r_46[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_92 = result_reg_r_46[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_93 = result_reg_r_46[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_94 = result_reg_r_46[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_95 = result_reg_r_46[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_96 = result_reg_r_46[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_97 = result_reg_r_46[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_98 = result_reg_r_46[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_99 = result_reg_r_46[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_100 = result_reg_r_46[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_101 = result_reg_r_46[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_102 = result_reg_r_46[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_103 = result_reg_r_46[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_104 = result_reg_r_46[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_93_105 = result_reg_r_46[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_47_hi_hi_hi_lo = {wire_res_93_98,wire_res_93_97,wire_res_93_96,wire_res_93_95,wire_res_93_94,
    wire_res_93_93,wire_res_93_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_47_hi_hi_lo_lo = {wire_res_93_84,wire_res_93_83,wire_res_93_82,wire_res_93_81,wire_res_93_80,
    wire_res_93_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_47_hi_hi_lo = {wire_res_93_91,wire_res_93_90,wire_res_93_89,wire_res_93_88,wire_res_93_87,
    wire_res_93_86,wire_res_93_85,result_reg_w_47_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_47_hi_lo_hi_lo = {wire_res_93_71,wire_res_93_70,wire_res_93_69,wire_res_93_68,wire_res_93_67,
    wire_res_93_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_47_hi_lo_lo_lo = {wire_res_93_58,wire_res_93_57,wire_res_93_56,wire_res_93_55,wire_res_93_54,
    wire_res_93_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_47_hi_lo_lo = {wire_res_93_65,wire_res_93_64,wire_res_93_63,wire_res_93_62,wire_res_93_61,
    wire_res_93_60,wire_res_93_59,result_reg_w_47_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_47_hi_lo = {wire_res_93_78,wire_res_93_77,wire_res_93_76,wire_res_93_75,wire_res_93_74,
    wire_res_93_73,wire_res_93_72,result_reg_w_47_hi_lo_hi_lo,result_reg_w_47_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_47_hi = {wire_res_93_105,wire_res_93_104,wire_res_93_103,wire_res_93_102,wire_res_93_101,
    wire_res_93_100,wire_res_93_99,result_reg_w_47_hi_hi_hi_lo,result_reg_w_47_hi_hi_lo,result_reg_w_47_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_47_lo_hi_hi_lo = {wire_res_93_45,wire_res_93_44,wire_res_93_43,wire_res_93_42,wire_res_93_41,
    wire_res_93_40,wire_res_93_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_47_lo_hi_lo_lo = {wire_res_93_31,wire_res_93_30,wire_res_93_29,wire_res_93_28,wire_res_93_27,
    wire_res_93_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_47_lo_hi_lo = {wire_res_93_38,wire_res_93_37,wire_res_93_36,wire_res_93_35,wire_res_93_34,
    wire_res_93_33,wire_res_93_32,result_reg_w_47_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_47_lo_lo_hi_lo = {wire_res_93_18,wire_res_93_17,wire_res_93_16,wire_res_93_15,wire_res_93_14,
    wire_res_93_13}; // @[BinaryDesigns2.scala 231:46]
  wire [116:0] _T_11424 = {b_aux_reg_r_46, 11'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [116:0] _GEN_1318 = {{11'd0}, a_aux_reg_r_46}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_93_11 = _GEN_1318 >= _T_11424; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_47_lo_lo_lo_lo = {wire_res_93_5,wire_res_93_4,wire_res_93_3,wire_res_93_2,wire_res_93_1,
    wire_res_93_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_47_lo_lo_lo = {wire_res_93_12,wire_res_93_11,wire_res_93_10,wire_res_93_9,wire_res_93_8,
    wire_res_93_7,wire_res_93_6,result_reg_w_47_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_47_lo_lo = {wire_res_93_25,wire_res_93_24,wire_res_93_23,wire_res_93_22,wire_res_93_21,
    wire_res_93_20,wire_res_93_19,result_reg_w_47_lo_lo_hi_lo,result_reg_w_47_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_47_lo = {wire_res_93_52,wire_res_93_51,wire_res_93_50,wire_res_93_49,wire_res_93_48,
    wire_res_93_47,wire_res_93_46,result_reg_w_47_lo_hi_hi_lo,result_reg_w_47_lo_hi_lo,result_reg_w_47_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_47 = {result_reg_w_47_hi,result_reg_w_47_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_94_0 = result_reg_w_47[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_1 = result_reg_w_47[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_2 = result_reg_w_47[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_3 = result_reg_w_47[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_4 = result_reg_w_47[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_5 = result_reg_w_47[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_6 = result_reg_w_47[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_7 = result_reg_w_47[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_8 = result_reg_w_47[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_9 = result_reg_w_47[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_11 = result_reg_w_47[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_12 = result_reg_w_47[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_13 = result_reg_w_47[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_14 = result_reg_w_47[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_15 = result_reg_w_47[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_16 = result_reg_w_47[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_17 = result_reg_w_47[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_18 = result_reg_w_47[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_19 = result_reg_w_47[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_20 = result_reg_w_47[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_21 = result_reg_w_47[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_22 = result_reg_w_47[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_23 = result_reg_w_47[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_24 = result_reg_w_47[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_25 = result_reg_w_47[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_26 = result_reg_w_47[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_27 = result_reg_w_47[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_28 = result_reg_w_47[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_29 = result_reg_w_47[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_30 = result_reg_w_47[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_31 = result_reg_w_47[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_32 = result_reg_w_47[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_33 = result_reg_w_47[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_34 = result_reg_w_47[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_35 = result_reg_w_47[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_36 = result_reg_w_47[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_37 = result_reg_w_47[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_38 = result_reg_w_47[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_39 = result_reg_w_47[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_40 = result_reg_w_47[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_41 = result_reg_w_47[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_42 = result_reg_w_47[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_43 = result_reg_w_47[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_44 = result_reg_w_47[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_45 = result_reg_w_47[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_46 = result_reg_w_47[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_47 = result_reg_w_47[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_48 = result_reg_w_47[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_49 = result_reg_w_47[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_50 = result_reg_w_47[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_51 = result_reg_w_47[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_52 = result_reg_w_47[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_53 = result_reg_w_47[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_54 = result_reg_w_47[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_55 = result_reg_w_47[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_56 = result_reg_w_47[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_57 = result_reg_w_47[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_58 = result_reg_w_47[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_59 = result_reg_w_47[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_60 = result_reg_w_47[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_61 = result_reg_w_47[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_62 = result_reg_w_47[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_63 = result_reg_w_47[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_64 = result_reg_w_47[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_65 = result_reg_w_47[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_66 = result_reg_w_47[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_67 = result_reg_w_47[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_68 = result_reg_w_47[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_69 = result_reg_w_47[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_70 = result_reg_w_47[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_71 = result_reg_w_47[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_72 = result_reg_w_47[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_73 = result_reg_w_47[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_74 = result_reg_w_47[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_75 = result_reg_w_47[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_76 = result_reg_w_47[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_77 = result_reg_w_47[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_78 = result_reg_w_47[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_79 = result_reg_w_47[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_80 = result_reg_w_47[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_81 = result_reg_w_47[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_82 = result_reg_w_47[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_83 = result_reg_w_47[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_84 = result_reg_w_47[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_85 = result_reg_w_47[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_86 = result_reg_w_47[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_87 = result_reg_w_47[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_88 = result_reg_w_47[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_89 = result_reg_w_47[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_90 = result_reg_w_47[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_91 = result_reg_w_47[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_92 = result_reg_w_47[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_93 = result_reg_w_47[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_94 = result_reg_w_47[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_95 = result_reg_w_47[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_96 = result_reg_w_47[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_97 = result_reg_w_47[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_98 = result_reg_w_47[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_99 = result_reg_w_47[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_100 = result_reg_w_47[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_101 = result_reg_w_47[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_102 = result_reg_w_47[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_103 = result_reg_w_47[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_104 = result_reg_w_47[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_94_105 = result_reg_w_47[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_0 = result_reg_r_47[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_1 = result_reg_r_47[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_2 = result_reg_r_47[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_3 = result_reg_r_47[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_4 = result_reg_r_47[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_5 = result_reg_r_47[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_6 = result_reg_r_47[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_7 = result_reg_r_47[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_8 = result_reg_r_47[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_10 = result_reg_r_47[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_11 = result_reg_r_47[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_12 = result_reg_r_47[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_13 = result_reg_r_47[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_14 = result_reg_r_47[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_15 = result_reg_r_47[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_16 = result_reg_r_47[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_17 = result_reg_r_47[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_18 = result_reg_r_47[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_19 = result_reg_r_47[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_20 = result_reg_r_47[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_21 = result_reg_r_47[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_22 = result_reg_r_47[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_23 = result_reg_r_47[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_24 = result_reg_r_47[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_25 = result_reg_r_47[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_26 = result_reg_r_47[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_27 = result_reg_r_47[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_28 = result_reg_r_47[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_29 = result_reg_r_47[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_30 = result_reg_r_47[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_31 = result_reg_r_47[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_32 = result_reg_r_47[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_33 = result_reg_r_47[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_34 = result_reg_r_47[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_35 = result_reg_r_47[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_36 = result_reg_r_47[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_37 = result_reg_r_47[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_38 = result_reg_r_47[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_39 = result_reg_r_47[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_40 = result_reg_r_47[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_41 = result_reg_r_47[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_42 = result_reg_r_47[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_43 = result_reg_r_47[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_44 = result_reg_r_47[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_45 = result_reg_r_47[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_46 = result_reg_r_47[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_47 = result_reg_r_47[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_48 = result_reg_r_47[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_49 = result_reg_r_47[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_50 = result_reg_r_47[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_51 = result_reg_r_47[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_52 = result_reg_r_47[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_53 = result_reg_r_47[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_54 = result_reg_r_47[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_55 = result_reg_r_47[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_56 = result_reg_r_47[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_57 = result_reg_r_47[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_58 = result_reg_r_47[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_59 = result_reg_r_47[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_60 = result_reg_r_47[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_61 = result_reg_r_47[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_62 = result_reg_r_47[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_63 = result_reg_r_47[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_64 = result_reg_r_47[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_65 = result_reg_r_47[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_66 = result_reg_r_47[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_67 = result_reg_r_47[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_68 = result_reg_r_47[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_69 = result_reg_r_47[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_70 = result_reg_r_47[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_71 = result_reg_r_47[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_72 = result_reg_r_47[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_73 = result_reg_r_47[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_74 = result_reg_r_47[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_75 = result_reg_r_47[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_76 = result_reg_r_47[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_77 = result_reg_r_47[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_78 = result_reg_r_47[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_79 = result_reg_r_47[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_80 = result_reg_r_47[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_81 = result_reg_r_47[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_82 = result_reg_r_47[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_83 = result_reg_r_47[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_84 = result_reg_r_47[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_85 = result_reg_r_47[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_86 = result_reg_r_47[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_87 = result_reg_r_47[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_88 = result_reg_r_47[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_89 = result_reg_r_47[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_90 = result_reg_r_47[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_91 = result_reg_r_47[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_92 = result_reg_r_47[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_93 = result_reg_r_47[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_94 = result_reg_r_47[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_95 = result_reg_r_47[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_96 = result_reg_r_47[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_97 = result_reg_r_47[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_98 = result_reg_r_47[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_99 = result_reg_r_47[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_100 = result_reg_r_47[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_101 = result_reg_r_47[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_102 = result_reg_r_47[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_103 = result_reg_r_47[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_104 = result_reg_r_47[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_95_105 = result_reg_r_47[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_48_hi_hi_hi_lo = {wire_res_95_98,wire_res_95_97,wire_res_95_96,wire_res_95_95,wire_res_95_94,
    wire_res_95_93,wire_res_95_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_48_hi_hi_lo_lo = {wire_res_95_84,wire_res_95_83,wire_res_95_82,wire_res_95_81,wire_res_95_80,
    wire_res_95_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_48_hi_hi_lo = {wire_res_95_91,wire_res_95_90,wire_res_95_89,wire_res_95_88,wire_res_95_87,
    wire_res_95_86,wire_res_95_85,result_reg_w_48_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_48_hi_lo_hi_lo = {wire_res_95_71,wire_res_95_70,wire_res_95_69,wire_res_95_68,wire_res_95_67,
    wire_res_95_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_48_hi_lo_lo_lo = {wire_res_95_58,wire_res_95_57,wire_res_95_56,wire_res_95_55,wire_res_95_54,
    wire_res_95_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_48_hi_lo_lo = {wire_res_95_65,wire_res_95_64,wire_res_95_63,wire_res_95_62,wire_res_95_61,
    wire_res_95_60,wire_res_95_59,result_reg_w_48_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_48_hi_lo = {wire_res_95_78,wire_res_95_77,wire_res_95_76,wire_res_95_75,wire_res_95_74,
    wire_res_95_73,wire_res_95_72,result_reg_w_48_hi_lo_hi_lo,result_reg_w_48_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_48_hi = {wire_res_95_105,wire_res_95_104,wire_res_95_103,wire_res_95_102,wire_res_95_101,
    wire_res_95_100,wire_res_95_99,result_reg_w_48_hi_hi_hi_lo,result_reg_w_48_hi_hi_lo,result_reg_w_48_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_48_lo_hi_hi_lo = {wire_res_95_45,wire_res_95_44,wire_res_95_43,wire_res_95_42,wire_res_95_41,
    wire_res_95_40,wire_res_95_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_48_lo_hi_lo_lo = {wire_res_95_31,wire_res_95_30,wire_res_95_29,wire_res_95_28,wire_res_95_27,
    wire_res_95_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_48_lo_hi_lo = {wire_res_95_38,wire_res_95_37,wire_res_95_36,wire_res_95_35,wire_res_95_34,
    wire_res_95_33,wire_res_95_32,result_reg_w_48_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_48_lo_lo_hi_lo = {wire_res_95_18,wire_res_95_17,wire_res_95_16,wire_res_95_15,wire_res_95_14,
    wire_res_95_13}; // @[BinaryDesigns2.scala 231:46]
  wire [114:0] _T_11428 = {b_aux_reg_r_47, 9'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [114:0] _GEN_1319 = {{9'd0}, a_aux_reg_r_47}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_95_9 = _GEN_1319 >= _T_11428; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_48_lo_lo_lo_lo = {wire_res_95_5,wire_res_95_4,wire_res_95_3,wire_res_95_2,wire_res_95_1,
    wire_res_95_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_48_lo_lo_lo = {wire_res_95_12,wire_res_95_11,wire_res_95_10,wire_res_95_9,wire_res_95_8,
    wire_res_95_7,wire_res_95_6,result_reg_w_48_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_48_lo_lo = {wire_res_95_25,wire_res_95_24,wire_res_95_23,wire_res_95_22,wire_res_95_21,
    wire_res_95_20,wire_res_95_19,result_reg_w_48_lo_lo_hi_lo,result_reg_w_48_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_48_lo = {wire_res_95_52,wire_res_95_51,wire_res_95_50,wire_res_95_49,wire_res_95_48,
    wire_res_95_47,wire_res_95_46,result_reg_w_48_lo_hi_hi_lo,result_reg_w_48_lo_hi_lo,result_reg_w_48_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_48 = {result_reg_w_48_hi,result_reg_w_48_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_96_0 = result_reg_w_48[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_1 = result_reg_w_48[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_2 = result_reg_w_48[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_3 = result_reg_w_48[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_4 = result_reg_w_48[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_5 = result_reg_w_48[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_6 = result_reg_w_48[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_7 = result_reg_w_48[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_9 = result_reg_w_48[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_10 = result_reg_w_48[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_11 = result_reg_w_48[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_12 = result_reg_w_48[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_13 = result_reg_w_48[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_14 = result_reg_w_48[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_15 = result_reg_w_48[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_16 = result_reg_w_48[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_17 = result_reg_w_48[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_18 = result_reg_w_48[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_19 = result_reg_w_48[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_20 = result_reg_w_48[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_21 = result_reg_w_48[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_22 = result_reg_w_48[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_23 = result_reg_w_48[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_24 = result_reg_w_48[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_25 = result_reg_w_48[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_26 = result_reg_w_48[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_27 = result_reg_w_48[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_28 = result_reg_w_48[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_29 = result_reg_w_48[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_30 = result_reg_w_48[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_31 = result_reg_w_48[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_32 = result_reg_w_48[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_33 = result_reg_w_48[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_34 = result_reg_w_48[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_35 = result_reg_w_48[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_36 = result_reg_w_48[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_37 = result_reg_w_48[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_38 = result_reg_w_48[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_39 = result_reg_w_48[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_40 = result_reg_w_48[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_41 = result_reg_w_48[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_42 = result_reg_w_48[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_43 = result_reg_w_48[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_44 = result_reg_w_48[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_45 = result_reg_w_48[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_46 = result_reg_w_48[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_47 = result_reg_w_48[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_48 = result_reg_w_48[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_49 = result_reg_w_48[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_50 = result_reg_w_48[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_51 = result_reg_w_48[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_52 = result_reg_w_48[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_53 = result_reg_w_48[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_54 = result_reg_w_48[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_55 = result_reg_w_48[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_56 = result_reg_w_48[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_57 = result_reg_w_48[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_58 = result_reg_w_48[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_59 = result_reg_w_48[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_60 = result_reg_w_48[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_61 = result_reg_w_48[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_62 = result_reg_w_48[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_63 = result_reg_w_48[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_64 = result_reg_w_48[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_65 = result_reg_w_48[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_66 = result_reg_w_48[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_67 = result_reg_w_48[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_68 = result_reg_w_48[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_69 = result_reg_w_48[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_70 = result_reg_w_48[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_71 = result_reg_w_48[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_72 = result_reg_w_48[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_73 = result_reg_w_48[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_74 = result_reg_w_48[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_75 = result_reg_w_48[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_76 = result_reg_w_48[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_77 = result_reg_w_48[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_78 = result_reg_w_48[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_79 = result_reg_w_48[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_80 = result_reg_w_48[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_81 = result_reg_w_48[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_82 = result_reg_w_48[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_83 = result_reg_w_48[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_84 = result_reg_w_48[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_85 = result_reg_w_48[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_86 = result_reg_w_48[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_87 = result_reg_w_48[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_88 = result_reg_w_48[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_89 = result_reg_w_48[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_90 = result_reg_w_48[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_91 = result_reg_w_48[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_92 = result_reg_w_48[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_93 = result_reg_w_48[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_94 = result_reg_w_48[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_95 = result_reg_w_48[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_96 = result_reg_w_48[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_97 = result_reg_w_48[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_98 = result_reg_w_48[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_99 = result_reg_w_48[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_100 = result_reg_w_48[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_101 = result_reg_w_48[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_102 = result_reg_w_48[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_103 = result_reg_w_48[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_104 = result_reg_w_48[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_96_105 = result_reg_w_48[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_0 = result_reg_r_48[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_1 = result_reg_r_48[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_2 = result_reg_r_48[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_3 = result_reg_r_48[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_4 = result_reg_r_48[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_5 = result_reg_r_48[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_6 = result_reg_r_48[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_8 = result_reg_r_48[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_9 = result_reg_r_48[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_10 = result_reg_r_48[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_11 = result_reg_r_48[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_12 = result_reg_r_48[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_13 = result_reg_r_48[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_14 = result_reg_r_48[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_15 = result_reg_r_48[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_16 = result_reg_r_48[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_17 = result_reg_r_48[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_18 = result_reg_r_48[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_19 = result_reg_r_48[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_20 = result_reg_r_48[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_21 = result_reg_r_48[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_22 = result_reg_r_48[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_23 = result_reg_r_48[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_24 = result_reg_r_48[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_25 = result_reg_r_48[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_26 = result_reg_r_48[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_27 = result_reg_r_48[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_28 = result_reg_r_48[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_29 = result_reg_r_48[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_30 = result_reg_r_48[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_31 = result_reg_r_48[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_32 = result_reg_r_48[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_33 = result_reg_r_48[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_34 = result_reg_r_48[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_35 = result_reg_r_48[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_36 = result_reg_r_48[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_37 = result_reg_r_48[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_38 = result_reg_r_48[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_39 = result_reg_r_48[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_40 = result_reg_r_48[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_41 = result_reg_r_48[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_42 = result_reg_r_48[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_43 = result_reg_r_48[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_44 = result_reg_r_48[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_45 = result_reg_r_48[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_46 = result_reg_r_48[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_47 = result_reg_r_48[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_48 = result_reg_r_48[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_49 = result_reg_r_48[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_50 = result_reg_r_48[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_51 = result_reg_r_48[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_52 = result_reg_r_48[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_53 = result_reg_r_48[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_54 = result_reg_r_48[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_55 = result_reg_r_48[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_56 = result_reg_r_48[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_57 = result_reg_r_48[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_58 = result_reg_r_48[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_59 = result_reg_r_48[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_60 = result_reg_r_48[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_61 = result_reg_r_48[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_62 = result_reg_r_48[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_63 = result_reg_r_48[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_64 = result_reg_r_48[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_65 = result_reg_r_48[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_66 = result_reg_r_48[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_67 = result_reg_r_48[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_68 = result_reg_r_48[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_69 = result_reg_r_48[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_70 = result_reg_r_48[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_71 = result_reg_r_48[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_72 = result_reg_r_48[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_73 = result_reg_r_48[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_74 = result_reg_r_48[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_75 = result_reg_r_48[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_76 = result_reg_r_48[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_77 = result_reg_r_48[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_78 = result_reg_r_48[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_79 = result_reg_r_48[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_80 = result_reg_r_48[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_81 = result_reg_r_48[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_82 = result_reg_r_48[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_83 = result_reg_r_48[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_84 = result_reg_r_48[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_85 = result_reg_r_48[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_86 = result_reg_r_48[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_87 = result_reg_r_48[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_88 = result_reg_r_48[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_89 = result_reg_r_48[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_90 = result_reg_r_48[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_91 = result_reg_r_48[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_92 = result_reg_r_48[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_93 = result_reg_r_48[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_94 = result_reg_r_48[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_95 = result_reg_r_48[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_96 = result_reg_r_48[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_97 = result_reg_r_48[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_98 = result_reg_r_48[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_99 = result_reg_r_48[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_100 = result_reg_r_48[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_101 = result_reg_r_48[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_102 = result_reg_r_48[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_103 = result_reg_r_48[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_104 = result_reg_r_48[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_97_105 = result_reg_r_48[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_49_hi_hi_hi_lo = {wire_res_97_98,wire_res_97_97,wire_res_97_96,wire_res_97_95,wire_res_97_94,
    wire_res_97_93,wire_res_97_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_49_hi_hi_lo_lo = {wire_res_97_84,wire_res_97_83,wire_res_97_82,wire_res_97_81,wire_res_97_80,
    wire_res_97_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_49_hi_hi_lo = {wire_res_97_91,wire_res_97_90,wire_res_97_89,wire_res_97_88,wire_res_97_87,
    wire_res_97_86,wire_res_97_85,result_reg_w_49_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_49_hi_lo_hi_lo = {wire_res_97_71,wire_res_97_70,wire_res_97_69,wire_res_97_68,wire_res_97_67,
    wire_res_97_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_49_hi_lo_lo_lo = {wire_res_97_58,wire_res_97_57,wire_res_97_56,wire_res_97_55,wire_res_97_54,
    wire_res_97_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_49_hi_lo_lo = {wire_res_97_65,wire_res_97_64,wire_res_97_63,wire_res_97_62,wire_res_97_61,
    wire_res_97_60,wire_res_97_59,result_reg_w_49_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_49_hi_lo = {wire_res_97_78,wire_res_97_77,wire_res_97_76,wire_res_97_75,wire_res_97_74,
    wire_res_97_73,wire_res_97_72,result_reg_w_49_hi_lo_hi_lo,result_reg_w_49_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_49_hi = {wire_res_97_105,wire_res_97_104,wire_res_97_103,wire_res_97_102,wire_res_97_101,
    wire_res_97_100,wire_res_97_99,result_reg_w_49_hi_hi_hi_lo,result_reg_w_49_hi_hi_lo,result_reg_w_49_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_49_lo_hi_hi_lo = {wire_res_97_45,wire_res_97_44,wire_res_97_43,wire_res_97_42,wire_res_97_41,
    wire_res_97_40,wire_res_97_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_49_lo_hi_lo_lo = {wire_res_97_31,wire_res_97_30,wire_res_97_29,wire_res_97_28,wire_res_97_27,
    wire_res_97_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_49_lo_hi_lo = {wire_res_97_38,wire_res_97_37,wire_res_97_36,wire_res_97_35,wire_res_97_34,
    wire_res_97_33,wire_res_97_32,result_reg_w_49_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_49_lo_lo_hi_lo = {wire_res_97_18,wire_res_97_17,wire_res_97_16,wire_res_97_15,wire_res_97_14,
    wire_res_97_13}; // @[BinaryDesigns2.scala 231:46]
  wire [112:0] _T_11432 = {b_aux_reg_r_48, 7'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [112:0] _GEN_1320 = {{7'd0}, a_aux_reg_r_48}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_97_7 = _GEN_1320 >= _T_11432; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_49_lo_lo_lo_lo = {wire_res_97_5,wire_res_97_4,wire_res_97_3,wire_res_97_2,wire_res_97_1,
    wire_res_97_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_49_lo_lo_lo = {wire_res_97_12,wire_res_97_11,wire_res_97_10,wire_res_97_9,wire_res_97_8,
    wire_res_97_7,wire_res_97_6,result_reg_w_49_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_49_lo_lo = {wire_res_97_25,wire_res_97_24,wire_res_97_23,wire_res_97_22,wire_res_97_21,
    wire_res_97_20,wire_res_97_19,result_reg_w_49_lo_lo_hi_lo,result_reg_w_49_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_49_lo = {wire_res_97_52,wire_res_97_51,wire_res_97_50,wire_res_97_49,wire_res_97_48,
    wire_res_97_47,wire_res_97_46,result_reg_w_49_lo_hi_hi_lo,result_reg_w_49_lo_hi_lo,result_reg_w_49_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_49 = {result_reg_w_49_hi,result_reg_w_49_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_98_0 = result_reg_w_49[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_1 = result_reg_w_49[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_2 = result_reg_w_49[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_3 = result_reg_w_49[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_4 = result_reg_w_49[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_5 = result_reg_w_49[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_7 = result_reg_w_49[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_8 = result_reg_w_49[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_9 = result_reg_w_49[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_10 = result_reg_w_49[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_11 = result_reg_w_49[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_12 = result_reg_w_49[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_13 = result_reg_w_49[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_14 = result_reg_w_49[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_15 = result_reg_w_49[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_16 = result_reg_w_49[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_17 = result_reg_w_49[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_18 = result_reg_w_49[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_19 = result_reg_w_49[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_20 = result_reg_w_49[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_21 = result_reg_w_49[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_22 = result_reg_w_49[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_23 = result_reg_w_49[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_24 = result_reg_w_49[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_25 = result_reg_w_49[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_26 = result_reg_w_49[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_27 = result_reg_w_49[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_28 = result_reg_w_49[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_29 = result_reg_w_49[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_30 = result_reg_w_49[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_31 = result_reg_w_49[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_32 = result_reg_w_49[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_33 = result_reg_w_49[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_34 = result_reg_w_49[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_35 = result_reg_w_49[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_36 = result_reg_w_49[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_37 = result_reg_w_49[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_38 = result_reg_w_49[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_39 = result_reg_w_49[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_40 = result_reg_w_49[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_41 = result_reg_w_49[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_42 = result_reg_w_49[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_43 = result_reg_w_49[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_44 = result_reg_w_49[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_45 = result_reg_w_49[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_46 = result_reg_w_49[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_47 = result_reg_w_49[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_48 = result_reg_w_49[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_49 = result_reg_w_49[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_50 = result_reg_w_49[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_51 = result_reg_w_49[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_52 = result_reg_w_49[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_53 = result_reg_w_49[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_54 = result_reg_w_49[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_55 = result_reg_w_49[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_56 = result_reg_w_49[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_57 = result_reg_w_49[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_58 = result_reg_w_49[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_59 = result_reg_w_49[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_60 = result_reg_w_49[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_61 = result_reg_w_49[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_62 = result_reg_w_49[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_63 = result_reg_w_49[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_64 = result_reg_w_49[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_65 = result_reg_w_49[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_66 = result_reg_w_49[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_67 = result_reg_w_49[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_68 = result_reg_w_49[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_69 = result_reg_w_49[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_70 = result_reg_w_49[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_71 = result_reg_w_49[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_72 = result_reg_w_49[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_73 = result_reg_w_49[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_74 = result_reg_w_49[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_75 = result_reg_w_49[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_76 = result_reg_w_49[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_77 = result_reg_w_49[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_78 = result_reg_w_49[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_79 = result_reg_w_49[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_80 = result_reg_w_49[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_81 = result_reg_w_49[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_82 = result_reg_w_49[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_83 = result_reg_w_49[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_84 = result_reg_w_49[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_85 = result_reg_w_49[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_86 = result_reg_w_49[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_87 = result_reg_w_49[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_88 = result_reg_w_49[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_89 = result_reg_w_49[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_90 = result_reg_w_49[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_91 = result_reg_w_49[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_92 = result_reg_w_49[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_93 = result_reg_w_49[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_94 = result_reg_w_49[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_95 = result_reg_w_49[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_96 = result_reg_w_49[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_97 = result_reg_w_49[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_98 = result_reg_w_49[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_99 = result_reg_w_49[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_100 = result_reg_w_49[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_101 = result_reg_w_49[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_102 = result_reg_w_49[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_103 = result_reg_w_49[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_104 = result_reg_w_49[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_98_105 = result_reg_w_49[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_0 = result_reg_r_49[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_1 = result_reg_r_49[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_2 = result_reg_r_49[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_3 = result_reg_r_49[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_4 = result_reg_r_49[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_6 = result_reg_r_49[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_7 = result_reg_r_49[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_8 = result_reg_r_49[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_9 = result_reg_r_49[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_10 = result_reg_r_49[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_11 = result_reg_r_49[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_12 = result_reg_r_49[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_13 = result_reg_r_49[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_14 = result_reg_r_49[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_15 = result_reg_r_49[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_16 = result_reg_r_49[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_17 = result_reg_r_49[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_18 = result_reg_r_49[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_19 = result_reg_r_49[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_20 = result_reg_r_49[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_21 = result_reg_r_49[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_22 = result_reg_r_49[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_23 = result_reg_r_49[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_24 = result_reg_r_49[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_25 = result_reg_r_49[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_26 = result_reg_r_49[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_27 = result_reg_r_49[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_28 = result_reg_r_49[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_29 = result_reg_r_49[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_30 = result_reg_r_49[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_31 = result_reg_r_49[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_32 = result_reg_r_49[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_33 = result_reg_r_49[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_34 = result_reg_r_49[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_35 = result_reg_r_49[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_36 = result_reg_r_49[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_37 = result_reg_r_49[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_38 = result_reg_r_49[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_39 = result_reg_r_49[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_40 = result_reg_r_49[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_41 = result_reg_r_49[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_42 = result_reg_r_49[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_43 = result_reg_r_49[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_44 = result_reg_r_49[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_45 = result_reg_r_49[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_46 = result_reg_r_49[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_47 = result_reg_r_49[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_48 = result_reg_r_49[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_49 = result_reg_r_49[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_50 = result_reg_r_49[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_51 = result_reg_r_49[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_52 = result_reg_r_49[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_53 = result_reg_r_49[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_54 = result_reg_r_49[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_55 = result_reg_r_49[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_56 = result_reg_r_49[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_57 = result_reg_r_49[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_58 = result_reg_r_49[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_59 = result_reg_r_49[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_60 = result_reg_r_49[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_61 = result_reg_r_49[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_62 = result_reg_r_49[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_63 = result_reg_r_49[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_64 = result_reg_r_49[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_65 = result_reg_r_49[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_66 = result_reg_r_49[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_67 = result_reg_r_49[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_68 = result_reg_r_49[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_69 = result_reg_r_49[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_70 = result_reg_r_49[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_71 = result_reg_r_49[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_72 = result_reg_r_49[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_73 = result_reg_r_49[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_74 = result_reg_r_49[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_75 = result_reg_r_49[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_76 = result_reg_r_49[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_77 = result_reg_r_49[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_78 = result_reg_r_49[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_79 = result_reg_r_49[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_80 = result_reg_r_49[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_81 = result_reg_r_49[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_82 = result_reg_r_49[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_83 = result_reg_r_49[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_84 = result_reg_r_49[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_85 = result_reg_r_49[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_86 = result_reg_r_49[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_87 = result_reg_r_49[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_88 = result_reg_r_49[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_89 = result_reg_r_49[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_90 = result_reg_r_49[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_91 = result_reg_r_49[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_92 = result_reg_r_49[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_93 = result_reg_r_49[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_94 = result_reg_r_49[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_95 = result_reg_r_49[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_96 = result_reg_r_49[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_97 = result_reg_r_49[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_98 = result_reg_r_49[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_99 = result_reg_r_49[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_100 = result_reg_r_49[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_101 = result_reg_r_49[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_102 = result_reg_r_49[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_103 = result_reg_r_49[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_104 = result_reg_r_49[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_99_105 = result_reg_r_49[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_50_hi_hi_hi_lo = {wire_res_99_98,wire_res_99_97,wire_res_99_96,wire_res_99_95,wire_res_99_94,
    wire_res_99_93,wire_res_99_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_50_hi_hi_lo_lo = {wire_res_99_84,wire_res_99_83,wire_res_99_82,wire_res_99_81,wire_res_99_80,
    wire_res_99_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_50_hi_hi_lo = {wire_res_99_91,wire_res_99_90,wire_res_99_89,wire_res_99_88,wire_res_99_87,
    wire_res_99_86,wire_res_99_85,result_reg_w_50_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_50_hi_lo_hi_lo = {wire_res_99_71,wire_res_99_70,wire_res_99_69,wire_res_99_68,wire_res_99_67,
    wire_res_99_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_50_hi_lo_lo_lo = {wire_res_99_58,wire_res_99_57,wire_res_99_56,wire_res_99_55,wire_res_99_54,
    wire_res_99_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_50_hi_lo_lo = {wire_res_99_65,wire_res_99_64,wire_res_99_63,wire_res_99_62,wire_res_99_61,
    wire_res_99_60,wire_res_99_59,result_reg_w_50_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_50_hi_lo = {wire_res_99_78,wire_res_99_77,wire_res_99_76,wire_res_99_75,wire_res_99_74,
    wire_res_99_73,wire_res_99_72,result_reg_w_50_hi_lo_hi_lo,result_reg_w_50_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_50_hi = {wire_res_99_105,wire_res_99_104,wire_res_99_103,wire_res_99_102,wire_res_99_101,
    wire_res_99_100,wire_res_99_99,result_reg_w_50_hi_hi_hi_lo,result_reg_w_50_hi_hi_lo,result_reg_w_50_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_50_lo_hi_hi_lo = {wire_res_99_45,wire_res_99_44,wire_res_99_43,wire_res_99_42,wire_res_99_41,
    wire_res_99_40,wire_res_99_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_50_lo_hi_lo_lo = {wire_res_99_31,wire_res_99_30,wire_res_99_29,wire_res_99_28,wire_res_99_27,
    wire_res_99_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_50_lo_hi_lo = {wire_res_99_38,wire_res_99_37,wire_res_99_36,wire_res_99_35,wire_res_99_34,
    wire_res_99_33,wire_res_99_32,result_reg_w_50_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_50_lo_lo_hi_lo = {wire_res_99_18,wire_res_99_17,wire_res_99_16,wire_res_99_15,wire_res_99_14,
    wire_res_99_13}; // @[BinaryDesigns2.scala 231:46]
  wire [110:0] _T_11436 = {b_aux_reg_r_49, 5'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [110:0] _GEN_1321 = {{5'd0}, a_aux_reg_r_49}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_99_5 = _GEN_1321 >= _T_11436; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_50_lo_lo_lo_lo = {wire_res_99_5,wire_res_99_4,wire_res_99_3,wire_res_99_2,wire_res_99_1,
    wire_res_99_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_50_lo_lo_lo = {wire_res_99_12,wire_res_99_11,wire_res_99_10,wire_res_99_9,wire_res_99_8,
    wire_res_99_7,wire_res_99_6,result_reg_w_50_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_50_lo_lo = {wire_res_99_25,wire_res_99_24,wire_res_99_23,wire_res_99_22,wire_res_99_21,
    wire_res_99_20,wire_res_99_19,result_reg_w_50_lo_lo_hi_lo,result_reg_w_50_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_50_lo = {wire_res_99_52,wire_res_99_51,wire_res_99_50,wire_res_99_49,wire_res_99_48,
    wire_res_99_47,wire_res_99_46,result_reg_w_50_lo_hi_hi_lo,result_reg_w_50_lo_hi_lo,result_reg_w_50_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_50 = {result_reg_w_50_hi,result_reg_w_50_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_100_0 = result_reg_w_50[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_1 = result_reg_w_50[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_2 = result_reg_w_50[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_3 = result_reg_w_50[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_5 = result_reg_w_50[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_6 = result_reg_w_50[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_7 = result_reg_w_50[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_8 = result_reg_w_50[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_9 = result_reg_w_50[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_10 = result_reg_w_50[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_11 = result_reg_w_50[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_12 = result_reg_w_50[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_13 = result_reg_w_50[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_14 = result_reg_w_50[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_15 = result_reg_w_50[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_16 = result_reg_w_50[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_17 = result_reg_w_50[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_18 = result_reg_w_50[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_19 = result_reg_w_50[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_20 = result_reg_w_50[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_21 = result_reg_w_50[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_22 = result_reg_w_50[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_23 = result_reg_w_50[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_24 = result_reg_w_50[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_25 = result_reg_w_50[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_26 = result_reg_w_50[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_27 = result_reg_w_50[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_28 = result_reg_w_50[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_29 = result_reg_w_50[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_30 = result_reg_w_50[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_31 = result_reg_w_50[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_32 = result_reg_w_50[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_33 = result_reg_w_50[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_34 = result_reg_w_50[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_35 = result_reg_w_50[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_36 = result_reg_w_50[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_37 = result_reg_w_50[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_38 = result_reg_w_50[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_39 = result_reg_w_50[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_40 = result_reg_w_50[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_41 = result_reg_w_50[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_42 = result_reg_w_50[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_43 = result_reg_w_50[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_44 = result_reg_w_50[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_45 = result_reg_w_50[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_46 = result_reg_w_50[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_47 = result_reg_w_50[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_48 = result_reg_w_50[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_49 = result_reg_w_50[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_50 = result_reg_w_50[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_51 = result_reg_w_50[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_52 = result_reg_w_50[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_53 = result_reg_w_50[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_54 = result_reg_w_50[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_55 = result_reg_w_50[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_56 = result_reg_w_50[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_57 = result_reg_w_50[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_58 = result_reg_w_50[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_59 = result_reg_w_50[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_60 = result_reg_w_50[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_61 = result_reg_w_50[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_62 = result_reg_w_50[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_63 = result_reg_w_50[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_64 = result_reg_w_50[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_65 = result_reg_w_50[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_66 = result_reg_w_50[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_67 = result_reg_w_50[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_68 = result_reg_w_50[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_69 = result_reg_w_50[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_70 = result_reg_w_50[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_71 = result_reg_w_50[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_72 = result_reg_w_50[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_73 = result_reg_w_50[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_74 = result_reg_w_50[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_75 = result_reg_w_50[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_76 = result_reg_w_50[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_77 = result_reg_w_50[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_78 = result_reg_w_50[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_79 = result_reg_w_50[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_80 = result_reg_w_50[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_81 = result_reg_w_50[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_82 = result_reg_w_50[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_83 = result_reg_w_50[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_84 = result_reg_w_50[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_85 = result_reg_w_50[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_86 = result_reg_w_50[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_87 = result_reg_w_50[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_88 = result_reg_w_50[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_89 = result_reg_w_50[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_90 = result_reg_w_50[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_91 = result_reg_w_50[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_92 = result_reg_w_50[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_93 = result_reg_w_50[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_94 = result_reg_w_50[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_95 = result_reg_w_50[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_96 = result_reg_w_50[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_97 = result_reg_w_50[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_98 = result_reg_w_50[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_99 = result_reg_w_50[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_100 = result_reg_w_50[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_101 = result_reg_w_50[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_102 = result_reg_w_50[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_103 = result_reg_w_50[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_104 = result_reg_w_50[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_100_105 = result_reg_w_50[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_0 = result_reg_r_50[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_1 = result_reg_r_50[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_2 = result_reg_r_50[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_4 = result_reg_r_50[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_5 = result_reg_r_50[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_6 = result_reg_r_50[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_7 = result_reg_r_50[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_8 = result_reg_r_50[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_9 = result_reg_r_50[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_10 = result_reg_r_50[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_11 = result_reg_r_50[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_12 = result_reg_r_50[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_13 = result_reg_r_50[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_14 = result_reg_r_50[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_15 = result_reg_r_50[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_16 = result_reg_r_50[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_17 = result_reg_r_50[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_18 = result_reg_r_50[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_19 = result_reg_r_50[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_20 = result_reg_r_50[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_21 = result_reg_r_50[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_22 = result_reg_r_50[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_23 = result_reg_r_50[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_24 = result_reg_r_50[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_25 = result_reg_r_50[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_26 = result_reg_r_50[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_27 = result_reg_r_50[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_28 = result_reg_r_50[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_29 = result_reg_r_50[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_30 = result_reg_r_50[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_31 = result_reg_r_50[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_32 = result_reg_r_50[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_33 = result_reg_r_50[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_34 = result_reg_r_50[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_35 = result_reg_r_50[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_36 = result_reg_r_50[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_37 = result_reg_r_50[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_38 = result_reg_r_50[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_39 = result_reg_r_50[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_40 = result_reg_r_50[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_41 = result_reg_r_50[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_42 = result_reg_r_50[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_43 = result_reg_r_50[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_44 = result_reg_r_50[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_45 = result_reg_r_50[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_46 = result_reg_r_50[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_47 = result_reg_r_50[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_48 = result_reg_r_50[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_49 = result_reg_r_50[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_50 = result_reg_r_50[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_51 = result_reg_r_50[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_52 = result_reg_r_50[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_53 = result_reg_r_50[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_54 = result_reg_r_50[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_55 = result_reg_r_50[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_56 = result_reg_r_50[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_57 = result_reg_r_50[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_58 = result_reg_r_50[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_59 = result_reg_r_50[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_60 = result_reg_r_50[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_61 = result_reg_r_50[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_62 = result_reg_r_50[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_63 = result_reg_r_50[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_64 = result_reg_r_50[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_65 = result_reg_r_50[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_66 = result_reg_r_50[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_67 = result_reg_r_50[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_68 = result_reg_r_50[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_69 = result_reg_r_50[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_70 = result_reg_r_50[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_71 = result_reg_r_50[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_72 = result_reg_r_50[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_73 = result_reg_r_50[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_74 = result_reg_r_50[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_75 = result_reg_r_50[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_76 = result_reg_r_50[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_77 = result_reg_r_50[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_78 = result_reg_r_50[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_79 = result_reg_r_50[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_80 = result_reg_r_50[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_81 = result_reg_r_50[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_82 = result_reg_r_50[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_83 = result_reg_r_50[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_84 = result_reg_r_50[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_85 = result_reg_r_50[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_86 = result_reg_r_50[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_87 = result_reg_r_50[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_88 = result_reg_r_50[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_89 = result_reg_r_50[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_90 = result_reg_r_50[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_91 = result_reg_r_50[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_92 = result_reg_r_50[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_93 = result_reg_r_50[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_94 = result_reg_r_50[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_95 = result_reg_r_50[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_96 = result_reg_r_50[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_97 = result_reg_r_50[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_98 = result_reg_r_50[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_99 = result_reg_r_50[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_100 = result_reg_r_50[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_101 = result_reg_r_50[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_102 = result_reg_r_50[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_103 = result_reg_r_50[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_104 = result_reg_r_50[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_101_105 = result_reg_r_50[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_51_hi_hi_hi_lo = {wire_res_101_98,wire_res_101_97,wire_res_101_96,wire_res_101_95,
    wire_res_101_94,wire_res_101_93,wire_res_101_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_51_hi_hi_lo_lo = {wire_res_101_84,wire_res_101_83,wire_res_101_82,wire_res_101_81,
    wire_res_101_80,wire_res_101_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_51_hi_hi_lo = {wire_res_101_91,wire_res_101_90,wire_res_101_89,wire_res_101_88,
    wire_res_101_87,wire_res_101_86,wire_res_101_85,result_reg_w_51_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_51_hi_lo_hi_lo = {wire_res_101_71,wire_res_101_70,wire_res_101_69,wire_res_101_68,
    wire_res_101_67,wire_res_101_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_51_hi_lo_lo_lo = {wire_res_101_58,wire_res_101_57,wire_res_101_56,wire_res_101_55,
    wire_res_101_54,wire_res_101_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_51_hi_lo_lo = {wire_res_101_65,wire_res_101_64,wire_res_101_63,wire_res_101_62,
    wire_res_101_61,wire_res_101_60,wire_res_101_59,result_reg_w_51_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_51_hi_lo = {wire_res_101_78,wire_res_101_77,wire_res_101_76,wire_res_101_75,wire_res_101_74,
    wire_res_101_73,wire_res_101_72,result_reg_w_51_hi_lo_hi_lo,result_reg_w_51_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_51_hi = {wire_res_101_105,wire_res_101_104,wire_res_101_103,wire_res_101_102,wire_res_101_101
    ,wire_res_101_100,wire_res_101_99,result_reg_w_51_hi_hi_hi_lo,result_reg_w_51_hi_hi_lo,result_reg_w_51_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_51_lo_hi_hi_lo = {wire_res_101_45,wire_res_101_44,wire_res_101_43,wire_res_101_42,
    wire_res_101_41,wire_res_101_40,wire_res_101_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_51_lo_hi_lo_lo = {wire_res_101_31,wire_res_101_30,wire_res_101_29,wire_res_101_28,
    wire_res_101_27,wire_res_101_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_51_lo_hi_lo = {wire_res_101_38,wire_res_101_37,wire_res_101_36,wire_res_101_35,
    wire_res_101_34,wire_res_101_33,wire_res_101_32,result_reg_w_51_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_51_lo_lo_hi_lo = {wire_res_101_18,wire_res_101_17,wire_res_101_16,wire_res_101_15,
    wire_res_101_14,wire_res_101_13}; // @[BinaryDesigns2.scala 231:46]
  wire [108:0] _T_11440 = {b_aux_reg_r_50, 3'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [108:0] _GEN_1322 = {{3'd0}, a_aux_reg_r_50}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_101_3 = _GEN_1322 >= _T_11440; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_51_lo_lo_lo_lo = {wire_res_101_5,wire_res_101_4,wire_res_101_3,wire_res_101_2,wire_res_101_1,
    wire_res_101_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_51_lo_lo_lo = {wire_res_101_12,wire_res_101_11,wire_res_101_10,wire_res_101_9,wire_res_101_8,
    wire_res_101_7,wire_res_101_6,result_reg_w_51_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_51_lo_lo = {wire_res_101_25,wire_res_101_24,wire_res_101_23,wire_res_101_22,wire_res_101_21,
    wire_res_101_20,wire_res_101_19,result_reg_w_51_lo_lo_hi_lo,result_reg_w_51_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_51_lo = {wire_res_101_52,wire_res_101_51,wire_res_101_50,wire_res_101_49,wire_res_101_48,
    wire_res_101_47,wire_res_101_46,result_reg_w_51_lo_hi_hi_lo,result_reg_w_51_lo_hi_lo,result_reg_w_51_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_51 = {result_reg_w_51_hi,result_reg_w_51_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_102_0 = result_reg_w_51[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_1 = result_reg_w_51[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_3 = result_reg_w_51[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_4 = result_reg_w_51[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_5 = result_reg_w_51[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_6 = result_reg_w_51[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_7 = result_reg_w_51[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_8 = result_reg_w_51[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_9 = result_reg_w_51[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_10 = result_reg_w_51[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_11 = result_reg_w_51[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_12 = result_reg_w_51[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_13 = result_reg_w_51[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_14 = result_reg_w_51[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_15 = result_reg_w_51[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_16 = result_reg_w_51[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_17 = result_reg_w_51[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_18 = result_reg_w_51[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_19 = result_reg_w_51[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_20 = result_reg_w_51[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_21 = result_reg_w_51[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_22 = result_reg_w_51[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_23 = result_reg_w_51[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_24 = result_reg_w_51[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_25 = result_reg_w_51[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_26 = result_reg_w_51[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_27 = result_reg_w_51[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_28 = result_reg_w_51[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_29 = result_reg_w_51[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_30 = result_reg_w_51[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_31 = result_reg_w_51[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_32 = result_reg_w_51[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_33 = result_reg_w_51[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_34 = result_reg_w_51[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_35 = result_reg_w_51[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_36 = result_reg_w_51[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_37 = result_reg_w_51[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_38 = result_reg_w_51[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_39 = result_reg_w_51[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_40 = result_reg_w_51[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_41 = result_reg_w_51[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_42 = result_reg_w_51[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_43 = result_reg_w_51[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_44 = result_reg_w_51[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_45 = result_reg_w_51[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_46 = result_reg_w_51[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_47 = result_reg_w_51[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_48 = result_reg_w_51[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_49 = result_reg_w_51[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_50 = result_reg_w_51[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_51 = result_reg_w_51[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_52 = result_reg_w_51[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_53 = result_reg_w_51[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_54 = result_reg_w_51[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_55 = result_reg_w_51[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_56 = result_reg_w_51[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_57 = result_reg_w_51[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_58 = result_reg_w_51[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_59 = result_reg_w_51[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_60 = result_reg_w_51[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_61 = result_reg_w_51[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_62 = result_reg_w_51[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_63 = result_reg_w_51[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_64 = result_reg_w_51[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_65 = result_reg_w_51[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_66 = result_reg_w_51[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_67 = result_reg_w_51[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_68 = result_reg_w_51[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_69 = result_reg_w_51[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_70 = result_reg_w_51[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_71 = result_reg_w_51[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_72 = result_reg_w_51[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_73 = result_reg_w_51[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_74 = result_reg_w_51[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_75 = result_reg_w_51[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_76 = result_reg_w_51[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_77 = result_reg_w_51[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_78 = result_reg_w_51[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_79 = result_reg_w_51[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_80 = result_reg_w_51[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_81 = result_reg_w_51[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_82 = result_reg_w_51[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_83 = result_reg_w_51[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_84 = result_reg_w_51[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_85 = result_reg_w_51[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_86 = result_reg_w_51[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_87 = result_reg_w_51[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_88 = result_reg_w_51[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_89 = result_reg_w_51[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_90 = result_reg_w_51[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_91 = result_reg_w_51[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_92 = result_reg_w_51[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_93 = result_reg_w_51[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_94 = result_reg_w_51[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_95 = result_reg_w_51[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_96 = result_reg_w_51[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_97 = result_reg_w_51[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_98 = result_reg_w_51[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_99 = result_reg_w_51[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_100 = result_reg_w_51[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_101 = result_reg_w_51[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_102 = result_reg_w_51[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_103 = result_reg_w_51[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_104 = result_reg_w_51[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_102_105 = result_reg_w_51[105]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_0 = result_reg_r_51[0]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_2 = result_reg_r_51[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_3 = result_reg_r_51[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_4 = result_reg_r_51[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_5 = result_reg_r_51[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_6 = result_reg_r_51[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_7 = result_reg_r_51[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_8 = result_reg_r_51[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_9 = result_reg_r_51[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_10 = result_reg_r_51[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_11 = result_reg_r_51[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_12 = result_reg_r_51[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_13 = result_reg_r_51[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_14 = result_reg_r_51[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_15 = result_reg_r_51[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_16 = result_reg_r_51[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_17 = result_reg_r_51[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_18 = result_reg_r_51[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_19 = result_reg_r_51[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_20 = result_reg_r_51[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_21 = result_reg_r_51[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_22 = result_reg_r_51[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_23 = result_reg_r_51[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_24 = result_reg_r_51[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_25 = result_reg_r_51[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_26 = result_reg_r_51[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_27 = result_reg_r_51[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_28 = result_reg_r_51[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_29 = result_reg_r_51[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_30 = result_reg_r_51[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_31 = result_reg_r_51[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_32 = result_reg_r_51[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_33 = result_reg_r_51[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_34 = result_reg_r_51[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_35 = result_reg_r_51[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_36 = result_reg_r_51[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_37 = result_reg_r_51[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_38 = result_reg_r_51[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_39 = result_reg_r_51[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_40 = result_reg_r_51[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_41 = result_reg_r_51[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_42 = result_reg_r_51[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_43 = result_reg_r_51[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_44 = result_reg_r_51[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_45 = result_reg_r_51[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_46 = result_reg_r_51[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_47 = result_reg_r_51[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_48 = result_reg_r_51[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_49 = result_reg_r_51[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_50 = result_reg_r_51[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_51 = result_reg_r_51[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_52 = result_reg_r_51[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_53 = result_reg_r_51[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_54 = result_reg_r_51[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_55 = result_reg_r_51[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_56 = result_reg_r_51[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_57 = result_reg_r_51[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_58 = result_reg_r_51[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_59 = result_reg_r_51[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_60 = result_reg_r_51[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_61 = result_reg_r_51[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_62 = result_reg_r_51[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_63 = result_reg_r_51[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_64 = result_reg_r_51[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_65 = result_reg_r_51[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_66 = result_reg_r_51[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_67 = result_reg_r_51[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_68 = result_reg_r_51[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_69 = result_reg_r_51[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_70 = result_reg_r_51[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_71 = result_reg_r_51[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_72 = result_reg_r_51[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_73 = result_reg_r_51[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_74 = result_reg_r_51[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_75 = result_reg_r_51[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_76 = result_reg_r_51[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_77 = result_reg_r_51[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_78 = result_reg_r_51[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_79 = result_reg_r_51[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_80 = result_reg_r_51[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_81 = result_reg_r_51[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_82 = result_reg_r_51[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_83 = result_reg_r_51[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_84 = result_reg_r_51[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_85 = result_reg_r_51[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_86 = result_reg_r_51[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_87 = result_reg_r_51[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_88 = result_reg_r_51[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_89 = result_reg_r_51[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_90 = result_reg_r_51[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_91 = result_reg_r_51[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_92 = result_reg_r_51[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_93 = result_reg_r_51[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_94 = result_reg_r_51[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_95 = result_reg_r_51[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_96 = result_reg_r_51[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_97 = result_reg_r_51[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_98 = result_reg_r_51[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_99 = result_reg_r_51[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_100 = result_reg_r_51[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_101 = result_reg_r_51[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_102 = result_reg_r_51[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_103 = result_reg_r_51[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_104 = result_reg_r_51[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_103_105 = result_reg_r_51[105]; // @[BinaryDesigns2.scala 192:62]
  wire [6:0] result_reg_w_52_hi_hi_hi_lo = {wire_res_103_98,wire_res_103_97,wire_res_103_96,wire_res_103_95,
    wire_res_103_94,wire_res_103_93,wire_res_103_92}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_52_hi_hi_lo_lo = {wire_res_103_84,wire_res_103_83,wire_res_103_82,wire_res_103_81,
    wire_res_103_80,wire_res_103_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_52_hi_hi_lo = {wire_res_103_91,wire_res_103_90,wire_res_103_89,wire_res_103_88,
    wire_res_103_87,wire_res_103_86,wire_res_103_85,result_reg_w_52_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_52_hi_lo_hi_lo = {wire_res_103_71,wire_res_103_70,wire_res_103_69,wire_res_103_68,
    wire_res_103_67,wire_res_103_66}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_52_hi_lo_lo_lo = {wire_res_103_58,wire_res_103_57,wire_res_103_56,wire_res_103_55,
    wire_res_103_54,wire_res_103_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_52_hi_lo_lo = {wire_res_103_65,wire_res_103_64,wire_res_103_63,wire_res_103_62,
    wire_res_103_61,wire_res_103_60,wire_res_103_59,result_reg_w_52_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_52_hi_lo = {wire_res_103_78,wire_res_103_77,wire_res_103_76,wire_res_103_75,wire_res_103_74,
    wire_res_103_73,wire_res_103_72,result_reg_w_52_hi_lo_hi_lo,result_reg_w_52_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_52_hi = {wire_res_103_105,wire_res_103_104,wire_res_103_103,wire_res_103_102,wire_res_103_101
    ,wire_res_103_100,wire_res_103_99,result_reg_w_52_hi_hi_hi_lo,result_reg_w_52_hi_hi_lo,result_reg_w_52_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_w_52_lo_hi_hi_lo = {wire_res_103_45,wire_res_103_44,wire_res_103_43,wire_res_103_42,
    wire_res_103_41,wire_res_103_40,wire_res_103_39}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_52_lo_hi_lo_lo = {wire_res_103_31,wire_res_103_30,wire_res_103_29,wire_res_103_28,
    wire_res_103_27,wire_res_103_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_52_lo_hi_lo = {wire_res_103_38,wire_res_103_37,wire_res_103_36,wire_res_103_35,
    wire_res_103_34,wire_res_103_33,wire_res_103_32,result_reg_w_52_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_w_52_lo_lo_hi_lo = {wire_res_103_18,wire_res_103_17,wire_res_103_16,wire_res_103_15,
    wire_res_103_14,wire_res_103_13}; // @[BinaryDesigns2.scala 231:46]
  wire [106:0] _T_11444 = {b_aux_reg_r_51, 1'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [106:0] _GEN_1323 = {{1'd0}, a_aux_reg_r_51}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_103_1 = _GEN_1323 >= _T_11444; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_w_52_lo_lo_lo_lo = {wire_res_103_5,wire_res_103_4,wire_res_103_3,wire_res_103_2,wire_res_103_1,
    wire_res_103_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_w_52_lo_lo_lo = {wire_res_103_12,wire_res_103_11,wire_res_103_10,wire_res_103_9,wire_res_103_8,
    wire_res_103_7,wire_res_103_6,result_reg_w_52_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_w_52_lo_lo = {wire_res_103_25,wire_res_103_24,wire_res_103_23,wire_res_103_22,wire_res_103_21,
    wire_res_103_20,wire_res_103_19,result_reg_w_52_lo_lo_hi_lo,result_reg_w_52_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_w_52_lo = {wire_res_103_52,wire_res_103_51,wire_res_103_50,wire_res_103_49,wire_res_103_48,
    wire_res_103_47,wire_res_103_46,result_reg_w_52_lo_hi_hi_lo,result_reg_w_52_lo_hi_lo,result_reg_w_52_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] result_reg_w_52 = {result_reg_w_52_hi,result_reg_w_52_lo}; // @[BinaryDesigns2.scala 231:46]
  wire  wire_res_104_1 = result_reg_w_52[1]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_2 = result_reg_w_52[2]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_3 = result_reg_w_52[3]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_4 = result_reg_w_52[4]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_5 = result_reg_w_52[5]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_6 = result_reg_w_52[6]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_7 = result_reg_w_52[7]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_8 = result_reg_w_52[8]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_9 = result_reg_w_52[9]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_10 = result_reg_w_52[10]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_11 = result_reg_w_52[11]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_12 = result_reg_w_52[12]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_13 = result_reg_w_52[13]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_14 = result_reg_w_52[14]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_15 = result_reg_w_52[15]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_16 = result_reg_w_52[16]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_17 = result_reg_w_52[17]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_18 = result_reg_w_52[18]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_19 = result_reg_w_52[19]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_20 = result_reg_w_52[20]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_21 = result_reg_w_52[21]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_22 = result_reg_w_52[22]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_23 = result_reg_w_52[23]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_24 = result_reg_w_52[24]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_25 = result_reg_w_52[25]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_26 = result_reg_w_52[26]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_27 = result_reg_w_52[27]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_28 = result_reg_w_52[28]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_29 = result_reg_w_52[29]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_30 = result_reg_w_52[30]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_31 = result_reg_w_52[31]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_32 = result_reg_w_52[32]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_33 = result_reg_w_52[33]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_34 = result_reg_w_52[34]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_35 = result_reg_w_52[35]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_36 = result_reg_w_52[36]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_37 = result_reg_w_52[37]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_38 = result_reg_w_52[38]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_39 = result_reg_w_52[39]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_40 = result_reg_w_52[40]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_41 = result_reg_w_52[41]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_42 = result_reg_w_52[42]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_43 = result_reg_w_52[43]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_44 = result_reg_w_52[44]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_45 = result_reg_w_52[45]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_46 = result_reg_w_52[46]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_47 = result_reg_w_52[47]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_48 = result_reg_w_52[48]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_49 = result_reg_w_52[49]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_50 = result_reg_w_52[50]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_51 = result_reg_w_52[51]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_52 = result_reg_w_52[52]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_53 = result_reg_w_52[53]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_54 = result_reg_w_52[54]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_55 = result_reg_w_52[55]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_56 = result_reg_w_52[56]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_57 = result_reg_w_52[57]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_58 = result_reg_w_52[58]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_59 = result_reg_w_52[59]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_60 = result_reg_w_52[60]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_61 = result_reg_w_52[61]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_62 = result_reg_w_52[62]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_63 = result_reg_w_52[63]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_64 = result_reg_w_52[64]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_65 = result_reg_w_52[65]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_66 = result_reg_w_52[66]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_67 = result_reg_w_52[67]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_68 = result_reg_w_52[68]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_69 = result_reg_w_52[69]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_70 = result_reg_w_52[70]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_71 = result_reg_w_52[71]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_72 = result_reg_w_52[72]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_73 = result_reg_w_52[73]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_74 = result_reg_w_52[74]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_75 = result_reg_w_52[75]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_76 = result_reg_w_52[76]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_77 = result_reg_w_52[77]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_78 = result_reg_w_52[78]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_79 = result_reg_w_52[79]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_80 = result_reg_w_52[80]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_81 = result_reg_w_52[81]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_82 = result_reg_w_52[82]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_83 = result_reg_w_52[83]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_84 = result_reg_w_52[84]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_85 = result_reg_w_52[85]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_86 = result_reg_w_52[86]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_87 = result_reg_w_52[87]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_88 = result_reg_w_52[88]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_89 = result_reg_w_52[89]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_90 = result_reg_w_52[90]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_91 = result_reg_w_52[91]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_92 = result_reg_w_52[92]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_93 = result_reg_w_52[93]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_94 = result_reg_w_52[94]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_95 = result_reg_w_52[95]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_96 = result_reg_w_52[96]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_97 = result_reg_w_52[97]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_98 = result_reg_w_52[98]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_99 = result_reg_w_52[99]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_100 = result_reg_w_52[100]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_101 = result_reg_w_52[101]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_102 = result_reg_w_52[102]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_103 = result_reg_w_52[103]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_104 = result_reg_w_52[104]; // @[BinaryDesigns2.scala 192:62]
  wire  wire_res_104_105 = result_reg_w_52[105]; // @[BinaryDesigns2.scala 192:62]
  wire [210:0] _GEN_1324 = {{105'd0}, io_in_a}; // @[BinaryDesigns2.scala 211:39]
  wire [105:0] a_aux_reg_w_0 = _GEN_1324[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [209:0] _GEN_1325 = {{104'd0}, a_aux_reg_w_0}; // @[BinaryDesigns2.scala 225:48]
  wire [208:0] _a_aux_reg_w_1_T_2 = _GEN_1272 - _T_11240; // @[BinaryDesigns2.scala 225:48]
  wire [208:0] _GEN_4 = wire_res_1_103 ? _a_aux_reg_w_1_T_2 : {{103'd0}, a_aux_reg_r_0}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [207:0] _T_11242 = {b_aux_reg_r_0, 102'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_1 = _GEN_4[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [207:0] _GEN_1327 = {{102'd0}, a_aux_reg_w_1}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_2_102 = _GEN_1327 >= _T_11242; // @[BinaryDesigns2.scala 224:35]
  wire [207:0] _a_aux_reg_r_1_T_2 = _GEN_1327 - _T_11242; // @[BinaryDesigns2.scala 225:48]
  wire [207:0] _GEN_6 = wire_res_2_102 ? _a_aux_reg_r_1_T_2 : {{102'd0}, a_aux_reg_w_1}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_1_lo_lo_lo_lo = {wire_res_2_5,wire_res_2_4,wire_res_2_3,wire_res_2_2,wire_res_2_1,wire_res_2_0
    }; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_1_lo_lo_lo = {wire_res_2_12,wire_res_2_11,wire_res_2_10,wire_res_2_9,wire_res_2_8,
    wire_res_2_7,wire_res_2_6,result_reg_r_1_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_1_lo_lo_hi_lo = {wire_res_2_18,wire_res_2_17,wire_res_2_16,wire_res_2_15,wire_res_2_14,
    wire_res_2_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_1_lo_lo = {wire_res_2_25,wire_res_2_24,wire_res_2_23,wire_res_2_22,wire_res_2_21,
    wire_res_2_20,wire_res_2_19,result_reg_r_1_lo_lo_hi_lo,result_reg_r_1_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_1_lo_hi_lo_lo = {wire_res_2_31,wire_res_2_30,wire_res_2_29,wire_res_2_28,wire_res_2_27,
    wire_res_2_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_1_lo_hi_lo = {wire_res_2_38,wire_res_2_37,wire_res_2_36,wire_res_2_35,wire_res_2_34,
    wire_res_2_33,wire_res_2_32,result_reg_r_1_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_1_lo_hi_hi_lo = {wire_res_2_45,wire_res_2_44,wire_res_2_43,wire_res_2_42,wire_res_2_41,
    wire_res_2_40,wire_res_2_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_1_lo = {wire_res_2_52,wire_res_2_51,wire_res_2_50,wire_res_2_49,wire_res_2_48,wire_res_2_47,
    wire_res_2_46,result_reg_r_1_lo_hi_hi_lo,result_reg_r_1_lo_hi_lo,result_reg_r_1_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_1_hi_lo_lo_lo = {wire_res_2_58,wire_res_2_57,wire_res_2_56,wire_res_2_55,wire_res_2_54,
    wire_res_2_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_1_hi_lo_lo = {wire_res_2_65,wire_res_2_64,wire_res_2_63,wire_res_2_62,wire_res_2_61,
    wire_res_2_60,wire_res_2_59,result_reg_r_1_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_1_hi_lo_hi_lo = {wire_res_2_71,wire_res_2_70,wire_res_2_69,wire_res_2_68,wire_res_2_67,
    wire_res_2_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_1_hi_lo = {wire_res_2_78,wire_res_2_77,wire_res_2_76,wire_res_2_75,wire_res_2_74,
    wire_res_2_73,wire_res_2_72,result_reg_r_1_hi_lo_hi_lo,result_reg_r_1_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_1_hi_hi_lo_lo = {wire_res_2_84,wire_res_2_83,wire_res_2_82,wire_res_2_81,wire_res_2_80,
    wire_res_2_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_1_hi_hi_lo = {wire_res_2_91,wire_res_2_90,wire_res_2_89,wire_res_2_88,wire_res_2_87,
    wire_res_2_86,wire_res_2_85,result_reg_r_1_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_1_hi_hi_hi_lo = {wire_res_2_98,wire_res_2_97,wire_res_2_96,wire_res_2_95,wire_res_2_94,
    wire_res_2_93,wire_res_2_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_1_hi = {wire_res_2_105,wire_res_2_104,wire_res_2_103,wire_res_2_102,wire_res_2_101,
    wire_res_2_100,wire_res_2_99,result_reg_r_1_hi_hi_hi_lo,result_reg_r_1_hi_hi_lo,result_reg_r_1_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_1_T = {result_reg_r_1_hi,result_reg_r_1_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [206:0] _a_aux_reg_w_2_T_2 = _GEN_1273 - _T_11244; // @[BinaryDesigns2.scala 225:48]
  wire [206:0] _GEN_8 = wire_res_3_101 ? _a_aux_reg_w_2_T_2 : {{101'd0}, a_aux_reg_r_1}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [205:0] _T_11246 = {b_aux_reg_r_1, 100'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_2 = _GEN_8[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [205:0] _GEN_1330 = {{100'd0}, a_aux_reg_w_2}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_4_100 = _GEN_1330 >= _T_11246; // @[BinaryDesigns2.scala 224:35]
  wire [205:0] _a_aux_reg_r_2_T_2 = _GEN_1330 - _T_11246; // @[BinaryDesigns2.scala 225:48]
  wire [205:0] _GEN_10 = wire_res_4_100 ? _a_aux_reg_r_2_T_2 : {{100'd0}, a_aux_reg_w_2}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_2_lo_lo_lo_lo = {wire_res_4_5,wire_res_4_4,wire_res_4_3,wire_res_4_2,wire_res_4_1,wire_res_4_0
    }; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_2_lo_lo_lo = {wire_res_4_12,wire_res_4_11,wire_res_4_10,wire_res_4_9,wire_res_4_8,
    wire_res_4_7,wire_res_4_6,result_reg_r_2_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_2_lo_lo_hi_lo = {wire_res_4_18,wire_res_4_17,wire_res_4_16,wire_res_4_15,wire_res_4_14,
    wire_res_4_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_2_lo_lo = {wire_res_4_25,wire_res_4_24,wire_res_4_23,wire_res_4_22,wire_res_4_21,
    wire_res_4_20,wire_res_4_19,result_reg_r_2_lo_lo_hi_lo,result_reg_r_2_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_2_lo_hi_lo_lo = {wire_res_4_31,wire_res_4_30,wire_res_4_29,wire_res_4_28,wire_res_4_27,
    wire_res_4_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_2_lo_hi_lo = {wire_res_4_38,wire_res_4_37,wire_res_4_36,wire_res_4_35,wire_res_4_34,
    wire_res_4_33,wire_res_4_32,result_reg_r_2_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_2_lo_hi_hi_lo = {wire_res_4_45,wire_res_4_44,wire_res_4_43,wire_res_4_42,wire_res_4_41,
    wire_res_4_40,wire_res_4_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_2_lo = {wire_res_4_52,wire_res_4_51,wire_res_4_50,wire_res_4_49,wire_res_4_48,wire_res_4_47,
    wire_res_4_46,result_reg_r_2_lo_hi_hi_lo,result_reg_r_2_lo_hi_lo,result_reg_r_2_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_2_hi_lo_lo_lo = {wire_res_4_58,wire_res_4_57,wire_res_4_56,wire_res_4_55,wire_res_4_54,
    wire_res_4_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_2_hi_lo_lo = {wire_res_4_65,wire_res_4_64,wire_res_4_63,wire_res_4_62,wire_res_4_61,
    wire_res_4_60,wire_res_4_59,result_reg_r_2_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_2_hi_lo_hi_lo = {wire_res_4_71,wire_res_4_70,wire_res_4_69,wire_res_4_68,wire_res_4_67,
    wire_res_4_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_2_hi_lo = {wire_res_4_78,wire_res_4_77,wire_res_4_76,wire_res_4_75,wire_res_4_74,
    wire_res_4_73,wire_res_4_72,result_reg_r_2_hi_lo_hi_lo,result_reg_r_2_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_2_hi_hi_lo_lo = {wire_res_4_84,wire_res_4_83,wire_res_4_82,wire_res_4_81,wire_res_4_80,
    wire_res_4_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_2_hi_hi_lo = {wire_res_4_91,wire_res_4_90,wire_res_4_89,wire_res_4_88,wire_res_4_87,
    wire_res_4_86,wire_res_4_85,result_reg_r_2_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_2_hi_hi_hi_lo = {wire_res_4_98,wire_res_4_97,wire_res_4_96,wire_res_4_95,wire_res_4_94,
    wire_res_4_93,wire_res_4_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_2_hi = {wire_res_4_105,wire_res_4_104,wire_res_4_103,wire_res_4_102,wire_res_4_101,
    wire_res_4_100,wire_res_4_99,result_reg_r_2_hi_hi_hi_lo,result_reg_r_2_hi_hi_lo,result_reg_r_2_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_2_T = {result_reg_r_2_hi,result_reg_r_2_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [204:0] _a_aux_reg_w_3_T_2 = _GEN_1274 - _T_11248; // @[BinaryDesigns2.scala 225:48]
  wire [204:0] _GEN_12 = wire_res_5_99 ? _a_aux_reg_w_3_T_2 : {{99'd0}, a_aux_reg_r_2}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [203:0] _T_11250 = {b_aux_reg_r_2, 98'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_3 = _GEN_12[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [203:0] _GEN_1333 = {{98'd0}, a_aux_reg_w_3}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_6_98 = _GEN_1333 >= _T_11250; // @[BinaryDesigns2.scala 224:35]
  wire [203:0] _a_aux_reg_r_3_T_2 = _GEN_1333 - _T_11250; // @[BinaryDesigns2.scala 225:48]
  wire [203:0] _GEN_14 = wire_res_6_98 ? _a_aux_reg_r_3_T_2 : {{98'd0}, a_aux_reg_w_3}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_3_lo_lo_lo_lo = {wire_res_6_5,wire_res_6_4,wire_res_6_3,wire_res_6_2,wire_res_6_1,wire_res_6_0
    }; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_3_lo_lo_lo = {wire_res_6_12,wire_res_6_11,wire_res_6_10,wire_res_6_9,wire_res_6_8,
    wire_res_6_7,wire_res_6_6,result_reg_r_3_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_3_lo_lo_hi_lo = {wire_res_6_18,wire_res_6_17,wire_res_6_16,wire_res_6_15,wire_res_6_14,
    wire_res_6_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_3_lo_lo = {wire_res_6_25,wire_res_6_24,wire_res_6_23,wire_res_6_22,wire_res_6_21,
    wire_res_6_20,wire_res_6_19,result_reg_r_3_lo_lo_hi_lo,result_reg_r_3_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_3_lo_hi_lo_lo = {wire_res_6_31,wire_res_6_30,wire_res_6_29,wire_res_6_28,wire_res_6_27,
    wire_res_6_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_3_lo_hi_lo = {wire_res_6_38,wire_res_6_37,wire_res_6_36,wire_res_6_35,wire_res_6_34,
    wire_res_6_33,wire_res_6_32,result_reg_r_3_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_3_lo_hi_hi_lo = {wire_res_6_45,wire_res_6_44,wire_res_6_43,wire_res_6_42,wire_res_6_41,
    wire_res_6_40,wire_res_6_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_3_lo = {wire_res_6_52,wire_res_6_51,wire_res_6_50,wire_res_6_49,wire_res_6_48,wire_res_6_47,
    wire_res_6_46,result_reg_r_3_lo_hi_hi_lo,result_reg_r_3_lo_hi_lo,result_reg_r_3_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_3_hi_lo_lo_lo = {wire_res_6_58,wire_res_6_57,wire_res_6_56,wire_res_6_55,wire_res_6_54,
    wire_res_6_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_3_hi_lo_lo = {wire_res_6_65,wire_res_6_64,wire_res_6_63,wire_res_6_62,wire_res_6_61,
    wire_res_6_60,wire_res_6_59,result_reg_r_3_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_3_hi_lo_hi_lo = {wire_res_6_71,wire_res_6_70,wire_res_6_69,wire_res_6_68,wire_res_6_67,
    wire_res_6_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_3_hi_lo = {wire_res_6_78,wire_res_6_77,wire_res_6_76,wire_res_6_75,wire_res_6_74,
    wire_res_6_73,wire_res_6_72,result_reg_r_3_hi_lo_hi_lo,result_reg_r_3_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_3_hi_hi_lo_lo = {wire_res_6_84,wire_res_6_83,wire_res_6_82,wire_res_6_81,wire_res_6_80,
    wire_res_6_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_3_hi_hi_lo = {wire_res_6_91,wire_res_6_90,wire_res_6_89,wire_res_6_88,wire_res_6_87,
    wire_res_6_86,wire_res_6_85,result_reg_r_3_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_3_hi_hi_hi_lo = {wire_res_6_98,wire_res_6_97,wire_res_6_96,wire_res_6_95,wire_res_6_94,
    wire_res_6_93,wire_res_6_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_3_hi = {wire_res_6_105,wire_res_6_104,wire_res_6_103,wire_res_6_102,wire_res_6_101,
    wire_res_6_100,wire_res_6_99,result_reg_r_3_hi_hi_hi_lo,result_reg_r_3_hi_hi_lo,result_reg_r_3_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_3_T = {result_reg_r_3_hi,result_reg_r_3_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [202:0] _a_aux_reg_w_4_T_2 = _GEN_1275 - _T_11252; // @[BinaryDesigns2.scala 225:48]
  wire [202:0] _GEN_16 = wire_res_7_97 ? _a_aux_reg_w_4_T_2 : {{97'd0}, a_aux_reg_r_3}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [201:0] _T_11254 = {b_aux_reg_r_3, 96'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_4 = _GEN_16[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [201:0] _GEN_1336 = {{96'd0}, a_aux_reg_w_4}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_8_96 = _GEN_1336 >= _T_11254; // @[BinaryDesigns2.scala 224:35]
  wire [201:0] _a_aux_reg_r_4_T_2 = _GEN_1336 - _T_11254; // @[BinaryDesigns2.scala 225:48]
  wire [201:0] _GEN_18 = wire_res_8_96 ? _a_aux_reg_r_4_T_2 : {{96'd0}, a_aux_reg_w_4}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_4_lo_lo_lo_lo = {wire_res_8_5,wire_res_8_4,wire_res_8_3,wire_res_8_2,wire_res_8_1,wire_res_8_0
    }; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_4_lo_lo_lo = {wire_res_8_12,wire_res_8_11,wire_res_8_10,wire_res_8_9,wire_res_8_8,
    wire_res_8_7,wire_res_8_6,result_reg_r_4_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_4_lo_lo_hi_lo = {wire_res_8_18,wire_res_8_17,wire_res_8_16,wire_res_8_15,wire_res_8_14,
    wire_res_8_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_4_lo_lo = {wire_res_8_25,wire_res_8_24,wire_res_8_23,wire_res_8_22,wire_res_8_21,
    wire_res_8_20,wire_res_8_19,result_reg_r_4_lo_lo_hi_lo,result_reg_r_4_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_4_lo_hi_lo_lo = {wire_res_8_31,wire_res_8_30,wire_res_8_29,wire_res_8_28,wire_res_8_27,
    wire_res_8_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_4_lo_hi_lo = {wire_res_8_38,wire_res_8_37,wire_res_8_36,wire_res_8_35,wire_res_8_34,
    wire_res_8_33,wire_res_8_32,result_reg_r_4_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_4_lo_hi_hi_lo = {wire_res_8_45,wire_res_8_44,wire_res_8_43,wire_res_8_42,wire_res_8_41,
    wire_res_8_40,wire_res_8_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_4_lo = {wire_res_8_52,wire_res_8_51,wire_res_8_50,wire_res_8_49,wire_res_8_48,wire_res_8_47,
    wire_res_8_46,result_reg_r_4_lo_hi_hi_lo,result_reg_r_4_lo_hi_lo,result_reg_r_4_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_4_hi_lo_lo_lo = {wire_res_8_58,wire_res_8_57,wire_res_8_56,wire_res_8_55,wire_res_8_54,
    wire_res_8_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_4_hi_lo_lo = {wire_res_8_65,wire_res_8_64,wire_res_8_63,wire_res_8_62,wire_res_8_61,
    wire_res_8_60,wire_res_8_59,result_reg_r_4_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_4_hi_lo_hi_lo = {wire_res_8_71,wire_res_8_70,wire_res_8_69,wire_res_8_68,wire_res_8_67,
    wire_res_8_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_4_hi_lo = {wire_res_8_78,wire_res_8_77,wire_res_8_76,wire_res_8_75,wire_res_8_74,
    wire_res_8_73,wire_res_8_72,result_reg_r_4_hi_lo_hi_lo,result_reg_r_4_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_4_hi_hi_lo_lo = {wire_res_8_84,wire_res_8_83,wire_res_8_82,wire_res_8_81,wire_res_8_80,
    wire_res_8_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_4_hi_hi_lo = {wire_res_8_91,wire_res_8_90,wire_res_8_89,wire_res_8_88,wire_res_8_87,
    wire_res_8_86,wire_res_8_85,result_reg_r_4_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_4_hi_hi_hi_lo = {wire_res_8_98,wire_res_8_97,wire_res_8_96,wire_res_8_95,wire_res_8_94,
    wire_res_8_93,wire_res_8_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_4_hi = {wire_res_8_105,wire_res_8_104,wire_res_8_103,wire_res_8_102,wire_res_8_101,
    wire_res_8_100,wire_res_8_99,result_reg_r_4_hi_hi_hi_lo,result_reg_r_4_hi_hi_lo,result_reg_r_4_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_4_T = {result_reg_r_4_hi,result_reg_r_4_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [200:0] _a_aux_reg_w_5_T_2 = _GEN_1276 - _T_11256; // @[BinaryDesigns2.scala 225:48]
  wire [200:0] _GEN_20 = wire_res_9_95 ? _a_aux_reg_w_5_T_2 : {{95'd0}, a_aux_reg_r_4}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [199:0] _T_11258 = {b_aux_reg_r_4, 94'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_5 = _GEN_20[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [199:0] _GEN_1339 = {{94'd0}, a_aux_reg_w_5}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_10_94 = _GEN_1339 >= _T_11258; // @[BinaryDesigns2.scala 224:35]
  wire [199:0] _a_aux_reg_r_5_T_2 = _GEN_1339 - _T_11258; // @[BinaryDesigns2.scala 225:48]
  wire [199:0] _GEN_22 = wire_res_10_94 ? _a_aux_reg_r_5_T_2 : {{94'd0}, a_aux_reg_w_5}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_5_lo_lo_lo_lo = {wire_res_10_5,wire_res_10_4,wire_res_10_3,wire_res_10_2,wire_res_10_1,
    wire_res_10_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_5_lo_lo_lo = {wire_res_10_12,wire_res_10_11,wire_res_10_10,wire_res_10_9,wire_res_10_8,
    wire_res_10_7,wire_res_10_6,result_reg_r_5_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_5_lo_lo_hi_lo = {wire_res_10_18,wire_res_10_17,wire_res_10_16,wire_res_10_15,wire_res_10_14,
    wire_res_10_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_5_lo_lo = {wire_res_10_25,wire_res_10_24,wire_res_10_23,wire_res_10_22,wire_res_10_21,
    wire_res_10_20,wire_res_10_19,result_reg_r_5_lo_lo_hi_lo,result_reg_r_5_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_5_lo_hi_lo_lo = {wire_res_10_31,wire_res_10_30,wire_res_10_29,wire_res_10_28,wire_res_10_27,
    wire_res_10_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_5_lo_hi_lo = {wire_res_10_38,wire_res_10_37,wire_res_10_36,wire_res_10_35,wire_res_10_34,
    wire_res_10_33,wire_res_10_32,result_reg_r_5_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_5_lo_hi_hi_lo = {wire_res_10_45,wire_res_10_44,wire_res_10_43,wire_res_10_42,wire_res_10_41,
    wire_res_10_40,wire_res_10_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_5_lo = {wire_res_10_52,wire_res_10_51,wire_res_10_50,wire_res_10_49,wire_res_10_48,
    wire_res_10_47,wire_res_10_46,result_reg_r_5_lo_hi_hi_lo,result_reg_r_5_lo_hi_lo,result_reg_r_5_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_5_hi_lo_lo_lo = {wire_res_10_58,wire_res_10_57,wire_res_10_56,wire_res_10_55,wire_res_10_54,
    wire_res_10_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_5_hi_lo_lo = {wire_res_10_65,wire_res_10_64,wire_res_10_63,wire_res_10_62,wire_res_10_61,
    wire_res_10_60,wire_res_10_59,result_reg_r_5_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_5_hi_lo_hi_lo = {wire_res_10_71,wire_res_10_70,wire_res_10_69,wire_res_10_68,wire_res_10_67,
    wire_res_10_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_5_hi_lo = {wire_res_10_78,wire_res_10_77,wire_res_10_76,wire_res_10_75,wire_res_10_74,
    wire_res_10_73,wire_res_10_72,result_reg_r_5_hi_lo_hi_lo,result_reg_r_5_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_5_hi_hi_lo_lo = {wire_res_10_84,wire_res_10_83,wire_res_10_82,wire_res_10_81,wire_res_10_80,
    wire_res_10_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_5_hi_hi_lo = {wire_res_10_91,wire_res_10_90,wire_res_10_89,wire_res_10_88,wire_res_10_87,
    wire_res_10_86,wire_res_10_85,result_reg_r_5_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_5_hi_hi_hi_lo = {wire_res_10_98,wire_res_10_97,wire_res_10_96,wire_res_10_95,wire_res_10_94,
    wire_res_10_93,wire_res_10_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_5_hi = {wire_res_10_105,wire_res_10_104,wire_res_10_103,wire_res_10_102,wire_res_10_101,
    wire_res_10_100,wire_res_10_99,result_reg_r_5_hi_hi_hi_lo,result_reg_r_5_hi_hi_lo,result_reg_r_5_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_5_T = {result_reg_r_5_hi,result_reg_r_5_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [198:0] _a_aux_reg_w_6_T_2 = _GEN_1277 - _T_11260; // @[BinaryDesigns2.scala 225:48]
  wire [198:0] _GEN_24 = wire_res_11_93 ? _a_aux_reg_w_6_T_2 : {{93'd0}, a_aux_reg_r_5}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [197:0] _T_11262 = {b_aux_reg_r_5, 92'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_6 = _GEN_24[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [197:0] _GEN_1342 = {{92'd0}, a_aux_reg_w_6}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_12_92 = _GEN_1342 >= _T_11262; // @[BinaryDesigns2.scala 224:35]
  wire [197:0] _a_aux_reg_r_6_T_2 = _GEN_1342 - _T_11262; // @[BinaryDesigns2.scala 225:48]
  wire [197:0] _GEN_26 = wire_res_12_92 ? _a_aux_reg_r_6_T_2 : {{92'd0}, a_aux_reg_w_6}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_6_lo_lo_lo_lo = {wire_res_12_5,wire_res_12_4,wire_res_12_3,wire_res_12_2,wire_res_12_1,
    wire_res_12_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_6_lo_lo_lo = {wire_res_12_12,wire_res_12_11,wire_res_12_10,wire_res_12_9,wire_res_12_8,
    wire_res_12_7,wire_res_12_6,result_reg_r_6_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_6_lo_lo_hi_lo = {wire_res_12_18,wire_res_12_17,wire_res_12_16,wire_res_12_15,wire_res_12_14,
    wire_res_12_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_6_lo_lo = {wire_res_12_25,wire_res_12_24,wire_res_12_23,wire_res_12_22,wire_res_12_21,
    wire_res_12_20,wire_res_12_19,result_reg_r_6_lo_lo_hi_lo,result_reg_r_6_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_6_lo_hi_lo_lo = {wire_res_12_31,wire_res_12_30,wire_res_12_29,wire_res_12_28,wire_res_12_27,
    wire_res_12_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_6_lo_hi_lo = {wire_res_12_38,wire_res_12_37,wire_res_12_36,wire_res_12_35,wire_res_12_34,
    wire_res_12_33,wire_res_12_32,result_reg_r_6_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_6_lo_hi_hi_lo = {wire_res_12_45,wire_res_12_44,wire_res_12_43,wire_res_12_42,wire_res_12_41,
    wire_res_12_40,wire_res_12_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_6_lo = {wire_res_12_52,wire_res_12_51,wire_res_12_50,wire_res_12_49,wire_res_12_48,
    wire_res_12_47,wire_res_12_46,result_reg_r_6_lo_hi_hi_lo,result_reg_r_6_lo_hi_lo,result_reg_r_6_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_6_hi_lo_lo_lo = {wire_res_12_58,wire_res_12_57,wire_res_12_56,wire_res_12_55,wire_res_12_54,
    wire_res_12_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_6_hi_lo_lo = {wire_res_12_65,wire_res_12_64,wire_res_12_63,wire_res_12_62,wire_res_12_61,
    wire_res_12_60,wire_res_12_59,result_reg_r_6_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_6_hi_lo_hi_lo = {wire_res_12_71,wire_res_12_70,wire_res_12_69,wire_res_12_68,wire_res_12_67,
    wire_res_12_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_6_hi_lo = {wire_res_12_78,wire_res_12_77,wire_res_12_76,wire_res_12_75,wire_res_12_74,
    wire_res_12_73,wire_res_12_72,result_reg_r_6_hi_lo_hi_lo,result_reg_r_6_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_6_hi_hi_lo_lo = {wire_res_12_84,wire_res_12_83,wire_res_12_82,wire_res_12_81,wire_res_12_80,
    wire_res_12_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_6_hi_hi_lo = {wire_res_12_91,wire_res_12_90,wire_res_12_89,wire_res_12_88,wire_res_12_87,
    wire_res_12_86,wire_res_12_85,result_reg_r_6_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_6_hi_hi_hi_lo = {wire_res_12_98,wire_res_12_97,wire_res_12_96,wire_res_12_95,wire_res_12_94,
    wire_res_12_93,wire_res_12_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_6_hi = {wire_res_12_105,wire_res_12_104,wire_res_12_103,wire_res_12_102,wire_res_12_101,
    wire_res_12_100,wire_res_12_99,result_reg_r_6_hi_hi_hi_lo,result_reg_r_6_hi_hi_lo,result_reg_r_6_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_6_T = {result_reg_r_6_hi,result_reg_r_6_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [196:0] _a_aux_reg_w_7_T_2 = _GEN_1278 - _T_11264; // @[BinaryDesigns2.scala 225:48]
  wire [196:0] _GEN_28 = wire_res_13_91 ? _a_aux_reg_w_7_T_2 : {{91'd0}, a_aux_reg_r_6}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [195:0] _T_11266 = {b_aux_reg_r_6, 90'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_7 = _GEN_28[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [195:0] _GEN_1345 = {{90'd0}, a_aux_reg_w_7}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_14_90 = _GEN_1345 >= _T_11266; // @[BinaryDesigns2.scala 224:35]
  wire [195:0] _a_aux_reg_r_7_T_2 = _GEN_1345 - _T_11266; // @[BinaryDesigns2.scala 225:48]
  wire [195:0] _GEN_30 = wire_res_14_90 ? _a_aux_reg_r_7_T_2 : {{90'd0}, a_aux_reg_w_7}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_7_lo_lo_lo_lo = {wire_res_14_5,wire_res_14_4,wire_res_14_3,wire_res_14_2,wire_res_14_1,
    wire_res_14_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_7_lo_lo_lo = {wire_res_14_12,wire_res_14_11,wire_res_14_10,wire_res_14_9,wire_res_14_8,
    wire_res_14_7,wire_res_14_6,result_reg_r_7_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_7_lo_lo_hi_lo = {wire_res_14_18,wire_res_14_17,wire_res_14_16,wire_res_14_15,wire_res_14_14,
    wire_res_14_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_7_lo_lo = {wire_res_14_25,wire_res_14_24,wire_res_14_23,wire_res_14_22,wire_res_14_21,
    wire_res_14_20,wire_res_14_19,result_reg_r_7_lo_lo_hi_lo,result_reg_r_7_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_7_lo_hi_lo_lo = {wire_res_14_31,wire_res_14_30,wire_res_14_29,wire_res_14_28,wire_res_14_27,
    wire_res_14_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_7_lo_hi_lo = {wire_res_14_38,wire_res_14_37,wire_res_14_36,wire_res_14_35,wire_res_14_34,
    wire_res_14_33,wire_res_14_32,result_reg_r_7_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_7_lo_hi_hi_lo = {wire_res_14_45,wire_res_14_44,wire_res_14_43,wire_res_14_42,wire_res_14_41,
    wire_res_14_40,wire_res_14_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_7_lo = {wire_res_14_52,wire_res_14_51,wire_res_14_50,wire_res_14_49,wire_res_14_48,
    wire_res_14_47,wire_res_14_46,result_reg_r_7_lo_hi_hi_lo,result_reg_r_7_lo_hi_lo,result_reg_r_7_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_7_hi_lo_lo_lo = {wire_res_14_58,wire_res_14_57,wire_res_14_56,wire_res_14_55,wire_res_14_54,
    wire_res_14_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_7_hi_lo_lo = {wire_res_14_65,wire_res_14_64,wire_res_14_63,wire_res_14_62,wire_res_14_61,
    wire_res_14_60,wire_res_14_59,result_reg_r_7_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_7_hi_lo_hi_lo = {wire_res_14_71,wire_res_14_70,wire_res_14_69,wire_res_14_68,wire_res_14_67,
    wire_res_14_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_7_hi_lo = {wire_res_14_78,wire_res_14_77,wire_res_14_76,wire_res_14_75,wire_res_14_74,
    wire_res_14_73,wire_res_14_72,result_reg_r_7_hi_lo_hi_lo,result_reg_r_7_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_7_hi_hi_lo_lo = {wire_res_14_84,wire_res_14_83,wire_res_14_82,wire_res_14_81,wire_res_14_80,
    wire_res_14_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_7_hi_hi_lo = {wire_res_14_91,wire_res_14_90,wire_res_14_89,wire_res_14_88,wire_res_14_87,
    wire_res_14_86,wire_res_14_85,result_reg_r_7_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_7_hi_hi_hi_lo = {wire_res_14_98,wire_res_14_97,wire_res_14_96,wire_res_14_95,wire_res_14_94,
    wire_res_14_93,wire_res_14_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_7_hi = {wire_res_14_105,wire_res_14_104,wire_res_14_103,wire_res_14_102,wire_res_14_101,
    wire_res_14_100,wire_res_14_99,result_reg_r_7_hi_hi_hi_lo,result_reg_r_7_hi_hi_lo,result_reg_r_7_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_7_T = {result_reg_r_7_hi,result_reg_r_7_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [194:0] _a_aux_reg_w_8_T_2 = _GEN_1279 - _T_11268; // @[BinaryDesigns2.scala 225:48]
  wire [194:0] _GEN_32 = wire_res_15_89 ? _a_aux_reg_w_8_T_2 : {{89'd0}, a_aux_reg_r_7}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [193:0] _T_11270 = {b_aux_reg_r_7, 88'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_8 = _GEN_32[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [193:0] _GEN_1348 = {{88'd0}, a_aux_reg_w_8}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_16_88 = _GEN_1348 >= _T_11270; // @[BinaryDesigns2.scala 224:35]
  wire [193:0] _a_aux_reg_r_8_T_2 = _GEN_1348 - _T_11270; // @[BinaryDesigns2.scala 225:48]
  wire [193:0] _GEN_34 = wire_res_16_88 ? _a_aux_reg_r_8_T_2 : {{88'd0}, a_aux_reg_w_8}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_8_lo_lo_lo_lo = {wire_res_16_5,wire_res_16_4,wire_res_16_3,wire_res_16_2,wire_res_16_1,
    wire_res_16_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_8_lo_lo_lo = {wire_res_16_12,wire_res_16_11,wire_res_16_10,wire_res_16_9,wire_res_16_8,
    wire_res_16_7,wire_res_16_6,result_reg_r_8_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_8_lo_lo_hi_lo = {wire_res_16_18,wire_res_16_17,wire_res_16_16,wire_res_16_15,wire_res_16_14,
    wire_res_16_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_8_lo_lo = {wire_res_16_25,wire_res_16_24,wire_res_16_23,wire_res_16_22,wire_res_16_21,
    wire_res_16_20,wire_res_16_19,result_reg_r_8_lo_lo_hi_lo,result_reg_r_8_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_8_lo_hi_lo_lo = {wire_res_16_31,wire_res_16_30,wire_res_16_29,wire_res_16_28,wire_res_16_27,
    wire_res_16_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_8_lo_hi_lo = {wire_res_16_38,wire_res_16_37,wire_res_16_36,wire_res_16_35,wire_res_16_34,
    wire_res_16_33,wire_res_16_32,result_reg_r_8_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_8_lo_hi_hi_lo = {wire_res_16_45,wire_res_16_44,wire_res_16_43,wire_res_16_42,wire_res_16_41,
    wire_res_16_40,wire_res_16_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_8_lo = {wire_res_16_52,wire_res_16_51,wire_res_16_50,wire_res_16_49,wire_res_16_48,
    wire_res_16_47,wire_res_16_46,result_reg_r_8_lo_hi_hi_lo,result_reg_r_8_lo_hi_lo,result_reg_r_8_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_8_hi_lo_lo_lo = {wire_res_16_58,wire_res_16_57,wire_res_16_56,wire_res_16_55,wire_res_16_54,
    wire_res_16_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_8_hi_lo_lo = {wire_res_16_65,wire_res_16_64,wire_res_16_63,wire_res_16_62,wire_res_16_61,
    wire_res_16_60,wire_res_16_59,result_reg_r_8_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_8_hi_lo_hi_lo = {wire_res_16_71,wire_res_16_70,wire_res_16_69,wire_res_16_68,wire_res_16_67,
    wire_res_16_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_8_hi_lo = {wire_res_16_78,wire_res_16_77,wire_res_16_76,wire_res_16_75,wire_res_16_74,
    wire_res_16_73,wire_res_16_72,result_reg_r_8_hi_lo_hi_lo,result_reg_r_8_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_8_hi_hi_lo_lo = {wire_res_16_84,wire_res_16_83,wire_res_16_82,wire_res_16_81,wire_res_16_80,
    wire_res_16_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_8_hi_hi_lo = {wire_res_16_91,wire_res_16_90,wire_res_16_89,wire_res_16_88,wire_res_16_87,
    wire_res_16_86,wire_res_16_85,result_reg_r_8_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_8_hi_hi_hi_lo = {wire_res_16_98,wire_res_16_97,wire_res_16_96,wire_res_16_95,wire_res_16_94,
    wire_res_16_93,wire_res_16_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_8_hi = {wire_res_16_105,wire_res_16_104,wire_res_16_103,wire_res_16_102,wire_res_16_101,
    wire_res_16_100,wire_res_16_99,result_reg_r_8_hi_hi_hi_lo,result_reg_r_8_hi_hi_lo,result_reg_r_8_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_8_T = {result_reg_r_8_hi,result_reg_r_8_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [192:0] _a_aux_reg_w_9_T_2 = _GEN_1280 - _T_11272; // @[BinaryDesigns2.scala 225:48]
  wire [192:0] _GEN_36 = wire_res_17_87 ? _a_aux_reg_w_9_T_2 : {{87'd0}, a_aux_reg_r_8}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [191:0] _T_11274 = {b_aux_reg_r_8, 86'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_9 = _GEN_36[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [191:0] _GEN_1351 = {{86'd0}, a_aux_reg_w_9}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_18_86 = _GEN_1351 >= _T_11274; // @[BinaryDesigns2.scala 224:35]
  wire [191:0] _a_aux_reg_r_9_T_2 = _GEN_1351 - _T_11274; // @[BinaryDesigns2.scala 225:48]
  wire [191:0] _GEN_38 = wire_res_18_86 ? _a_aux_reg_r_9_T_2 : {{86'd0}, a_aux_reg_w_9}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_9_lo_lo_lo_lo = {wire_res_18_5,wire_res_18_4,wire_res_18_3,wire_res_18_2,wire_res_18_1,
    wire_res_18_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_9_lo_lo_lo = {wire_res_18_12,wire_res_18_11,wire_res_18_10,wire_res_18_9,wire_res_18_8,
    wire_res_18_7,wire_res_18_6,result_reg_r_9_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_9_lo_lo_hi_lo = {wire_res_18_18,wire_res_18_17,wire_res_18_16,wire_res_18_15,wire_res_18_14,
    wire_res_18_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_9_lo_lo = {wire_res_18_25,wire_res_18_24,wire_res_18_23,wire_res_18_22,wire_res_18_21,
    wire_res_18_20,wire_res_18_19,result_reg_r_9_lo_lo_hi_lo,result_reg_r_9_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_9_lo_hi_lo_lo = {wire_res_18_31,wire_res_18_30,wire_res_18_29,wire_res_18_28,wire_res_18_27,
    wire_res_18_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_9_lo_hi_lo = {wire_res_18_38,wire_res_18_37,wire_res_18_36,wire_res_18_35,wire_res_18_34,
    wire_res_18_33,wire_res_18_32,result_reg_r_9_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_9_lo_hi_hi_lo = {wire_res_18_45,wire_res_18_44,wire_res_18_43,wire_res_18_42,wire_res_18_41,
    wire_res_18_40,wire_res_18_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_9_lo = {wire_res_18_52,wire_res_18_51,wire_res_18_50,wire_res_18_49,wire_res_18_48,
    wire_res_18_47,wire_res_18_46,result_reg_r_9_lo_hi_hi_lo,result_reg_r_9_lo_hi_lo,result_reg_r_9_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_9_hi_lo_lo_lo = {wire_res_18_58,wire_res_18_57,wire_res_18_56,wire_res_18_55,wire_res_18_54,
    wire_res_18_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_9_hi_lo_lo = {wire_res_18_65,wire_res_18_64,wire_res_18_63,wire_res_18_62,wire_res_18_61,
    wire_res_18_60,wire_res_18_59,result_reg_r_9_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_9_hi_lo_hi_lo = {wire_res_18_71,wire_res_18_70,wire_res_18_69,wire_res_18_68,wire_res_18_67,
    wire_res_18_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_9_hi_lo = {wire_res_18_78,wire_res_18_77,wire_res_18_76,wire_res_18_75,wire_res_18_74,
    wire_res_18_73,wire_res_18_72,result_reg_r_9_hi_lo_hi_lo,result_reg_r_9_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_9_hi_hi_lo_lo = {wire_res_18_84,wire_res_18_83,wire_res_18_82,wire_res_18_81,wire_res_18_80,
    wire_res_18_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_9_hi_hi_lo = {wire_res_18_91,wire_res_18_90,wire_res_18_89,wire_res_18_88,wire_res_18_87,
    wire_res_18_86,wire_res_18_85,result_reg_r_9_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_9_hi_hi_hi_lo = {wire_res_18_98,wire_res_18_97,wire_res_18_96,wire_res_18_95,wire_res_18_94,
    wire_res_18_93,wire_res_18_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_9_hi = {wire_res_18_105,wire_res_18_104,wire_res_18_103,wire_res_18_102,wire_res_18_101,
    wire_res_18_100,wire_res_18_99,result_reg_r_9_hi_hi_hi_lo,result_reg_r_9_hi_hi_lo,result_reg_r_9_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_9_T = {result_reg_r_9_hi,result_reg_r_9_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [190:0] _a_aux_reg_w_10_T_2 = _GEN_1281 - _T_11276; // @[BinaryDesigns2.scala 225:48]
  wire [190:0] _GEN_40 = wire_res_19_85 ? _a_aux_reg_w_10_T_2 : {{85'd0}, a_aux_reg_r_9}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [189:0] _T_11278 = {b_aux_reg_r_9, 84'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_10 = _GEN_40[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [189:0] _GEN_1354 = {{84'd0}, a_aux_reg_w_10}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_20_84 = _GEN_1354 >= _T_11278; // @[BinaryDesigns2.scala 224:35]
  wire [189:0] _a_aux_reg_r_10_T_2 = _GEN_1354 - _T_11278; // @[BinaryDesigns2.scala 225:48]
  wire [189:0] _GEN_42 = wire_res_20_84 ? _a_aux_reg_r_10_T_2 : {{84'd0}, a_aux_reg_w_10}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_10_lo_lo_lo_lo = {wire_res_20_5,wire_res_20_4,wire_res_20_3,wire_res_20_2,wire_res_20_1,
    wire_res_20_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_10_lo_lo_lo = {wire_res_20_12,wire_res_20_11,wire_res_20_10,wire_res_20_9,wire_res_20_8,
    wire_res_20_7,wire_res_20_6,result_reg_r_10_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_10_lo_lo_hi_lo = {wire_res_20_18,wire_res_20_17,wire_res_20_16,wire_res_20_15,wire_res_20_14,
    wire_res_20_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_10_lo_lo = {wire_res_20_25,wire_res_20_24,wire_res_20_23,wire_res_20_22,wire_res_20_21,
    wire_res_20_20,wire_res_20_19,result_reg_r_10_lo_lo_hi_lo,result_reg_r_10_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_10_lo_hi_lo_lo = {wire_res_20_31,wire_res_20_30,wire_res_20_29,wire_res_20_28,wire_res_20_27,
    wire_res_20_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_10_lo_hi_lo = {wire_res_20_38,wire_res_20_37,wire_res_20_36,wire_res_20_35,wire_res_20_34,
    wire_res_20_33,wire_res_20_32,result_reg_r_10_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_10_lo_hi_hi_lo = {wire_res_20_45,wire_res_20_44,wire_res_20_43,wire_res_20_42,wire_res_20_41,
    wire_res_20_40,wire_res_20_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_10_lo = {wire_res_20_52,wire_res_20_51,wire_res_20_50,wire_res_20_49,wire_res_20_48,
    wire_res_20_47,wire_res_20_46,result_reg_r_10_lo_hi_hi_lo,result_reg_r_10_lo_hi_lo,result_reg_r_10_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_10_hi_lo_lo_lo = {wire_res_20_58,wire_res_20_57,wire_res_20_56,wire_res_20_55,wire_res_20_54,
    wire_res_20_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_10_hi_lo_lo = {wire_res_20_65,wire_res_20_64,wire_res_20_63,wire_res_20_62,wire_res_20_61,
    wire_res_20_60,wire_res_20_59,result_reg_r_10_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_10_hi_lo_hi_lo = {wire_res_20_71,wire_res_20_70,wire_res_20_69,wire_res_20_68,wire_res_20_67,
    wire_res_20_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_10_hi_lo = {wire_res_20_78,wire_res_20_77,wire_res_20_76,wire_res_20_75,wire_res_20_74,
    wire_res_20_73,wire_res_20_72,result_reg_r_10_hi_lo_hi_lo,result_reg_r_10_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_10_hi_hi_lo_lo = {wire_res_20_84,wire_res_20_83,wire_res_20_82,wire_res_20_81,wire_res_20_80,
    wire_res_20_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_10_hi_hi_lo = {wire_res_20_91,wire_res_20_90,wire_res_20_89,wire_res_20_88,wire_res_20_87,
    wire_res_20_86,wire_res_20_85,result_reg_r_10_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_10_hi_hi_hi_lo = {wire_res_20_98,wire_res_20_97,wire_res_20_96,wire_res_20_95,wire_res_20_94,
    wire_res_20_93,wire_res_20_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_10_hi = {wire_res_20_105,wire_res_20_104,wire_res_20_103,wire_res_20_102,wire_res_20_101,
    wire_res_20_100,wire_res_20_99,result_reg_r_10_hi_hi_hi_lo,result_reg_r_10_hi_hi_lo,result_reg_r_10_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_10_T = {result_reg_r_10_hi,result_reg_r_10_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [188:0] _a_aux_reg_w_11_T_2 = _GEN_1282 - _T_11280; // @[BinaryDesigns2.scala 225:48]
  wire [188:0] _GEN_44 = wire_res_21_83 ? _a_aux_reg_w_11_T_2 : {{83'd0}, a_aux_reg_r_10}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [187:0] _T_11282 = {b_aux_reg_r_10, 82'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_11 = _GEN_44[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [187:0] _GEN_1357 = {{82'd0}, a_aux_reg_w_11}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_22_82 = _GEN_1357 >= _T_11282; // @[BinaryDesigns2.scala 224:35]
  wire [187:0] _a_aux_reg_r_11_T_2 = _GEN_1357 - _T_11282; // @[BinaryDesigns2.scala 225:48]
  wire [187:0] _GEN_46 = wire_res_22_82 ? _a_aux_reg_r_11_T_2 : {{82'd0}, a_aux_reg_w_11}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_11_lo_lo_lo_lo = {wire_res_22_5,wire_res_22_4,wire_res_22_3,wire_res_22_2,wire_res_22_1,
    wire_res_22_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_11_lo_lo_lo = {wire_res_22_12,wire_res_22_11,wire_res_22_10,wire_res_22_9,wire_res_22_8,
    wire_res_22_7,wire_res_22_6,result_reg_r_11_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_11_lo_lo_hi_lo = {wire_res_22_18,wire_res_22_17,wire_res_22_16,wire_res_22_15,wire_res_22_14,
    wire_res_22_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_11_lo_lo = {wire_res_22_25,wire_res_22_24,wire_res_22_23,wire_res_22_22,wire_res_22_21,
    wire_res_22_20,wire_res_22_19,result_reg_r_11_lo_lo_hi_lo,result_reg_r_11_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_11_lo_hi_lo_lo = {wire_res_22_31,wire_res_22_30,wire_res_22_29,wire_res_22_28,wire_res_22_27,
    wire_res_22_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_11_lo_hi_lo = {wire_res_22_38,wire_res_22_37,wire_res_22_36,wire_res_22_35,wire_res_22_34,
    wire_res_22_33,wire_res_22_32,result_reg_r_11_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_11_lo_hi_hi_lo = {wire_res_22_45,wire_res_22_44,wire_res_22_43,wire_res_22_42,wire_res_22_41,
    wire_res_22_40,wire_res_22_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_11_lo = {wire_res_22_52,wire_res_22_51,wire_res_22_50,wire_res_22_49,wire_res_22_48,
    wire_res_22_47,wire_res_22_46,result_reg_r_11_lo_hi_hi_lo,result_reg_r_11_lo_hi_lo,result_reg_r_11_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_11_hi_lo_lo_lo = {wire_res_22_58,wire_res_22_57,wire_res_22_56,wire_res_22_55,wire_res_22_54,
    wire_res_22_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_11_hi_lo_lo = {wire_res_22_65,wire_res_22_64,wire_res_22_63,wire_res_22_62,wire_res_22_61,
    wire_res_22_60,wire_res_22_59,result_reg_r_11_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_11_hi_lo_hi_lo = {wire_res_22_71,wire_res_22_70,wire_res_22_69,wire_res_22_68,wire_res_22_67,
    wire_res_22_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_11_hi_lo = {wire_res_22_78,wire_res_22_77,wire_res_22_76,wire_res_22_75,wire_res_22_74,
    wire_res_22_73,wire_res_22_72,result_reg_r_11_hi_lo_hi_lo,result_reg_r_11_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_11_hi_hi_lo_lo = {wire_res_22_84,wire_res_22_83,wire_res_22_82,wire_res_22_81,wire_res_22_80,
    wire_res_22_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_11_hi_hi_lo = {wire_res_22_91,wire_res_22_90,wire_res_22_89,wire_res_22_88,wire_res_22_87,
    wire_res_22_86,wire_res_22_85,result_reg_r_11_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_11_hi_hi_hi_lo = {wire_res_22_98,wire_res_22_97,wire_res_22_96,wire_res_22_95,wire_res_22_94,
    wire_res_22_93,wire_res_22_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_11_hi = {wire_res_22_105,wire_res_22_104,wire_res_22_103,wire_res_22_102,wire_res_22_101,
    wire_res_22_100,wire_res_22_99,result_reg_r_11_hi_hi_hi_lo,result_reg_r_11_hi_hi_lo,result_reg_r_11_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_11_T = {result_reg_r_11_hi,result_reg_r_11_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [186:0] _a_aux_reg_w_12_T_2 = _GEN_1283 - _T_11284; // @[BinaryDesigns2.scala 225:48]
  wire [186:0] _GEN_48 = wire_res_23_81 ? _a_aux_reg_w_12_T_2 : {{81'd0}, a_aux_reg_r_11}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [185:0] _T_11286 = {b_aux_reg_r_11, 80'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_12 = _GEN_48[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [185:0] _GEN_1360 = {{80'd0}, a_aux_reg_w_12}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_24_80 = _GEN_1360 >= _T_11286; // @[BinaryDesigns2.scala 224:35]
  wire [185:0] _a_aux_reg_r_12_T_2 = _GEN_1360 - _T_11286; // @[BinaryDesigns2.scala 225:48]
  wire [185:0] _GEN_50 = wire_res_24_80 ? _a_aux_reg_r_12_T_2 : {{80'd0}, a_aux_reg_w_12}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_12_lo_lo_lo_lo = {wire_res_24_5,wire_res_24_4,wire_res_24_3,wire_res_24_2,wire_res_24_1,
    wire_res_24_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_12_lo_lo_lo = {wire_res_24_12,wire_res_24_11,wire_res_24_10,wire_res_24_9,wire_res_24_8,
    wire_res_24_7,wire_res_24_6,result_reg_r_12_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_12_lo_lo_hi_lo = {wire_res_24_18,wire_res_24_17,wire_res_24_16,wire_res_24_15,wire_res_24_14,
    wire_res_24_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_12_lo_lo = {wire_res_24_25,wire_res_24_24,wire_res_24_23,wire_res_24_22,wire_res_24_21,
    wire_res_24_20,wire_res_24_19,result_reg_r_12_lo_lo_hi_lo,result_reg_r_12_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_12_lo_hi_lo_lo = {wire_res_24_31,wire_res_24_30,wire_res_24_29,wire_res_24_28,wire_res_24_27,
    wire_res_24_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_12_lo_hi_lo = {wire_res_24_38,wire_res_24_37,wire_res_24_36,wire_res_24_35,wire_res_24_34,
    wire_res_24_33,wire_res_24_32,result_reg_r_12_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_12_lo_hi_hi_lo = {wire_res_24_45,wire_res_24_44,wire_res_24_43,wire_res_24_42,wire_res_24_41,
    wire_res_24_40,wire_res_24_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_12_lo = {wire_res_24_52,wire_res_24_51,wire_res_24_50,wire_res_24_49,wire_res_24_48,
    wire_res_24_47,wire_res_24_46,result_reg_r_12_lo_hi_hi_lo,result_reg_r_12_lo_hi_lo,result_reg_r_12_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_12_hi_lo_lo_lo = {wire_res_24_58,wire_res_24_57,wire_res_24_56,wire_res_24_55,wire_res_24_54,
    wire_res_24_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_12_hi_lo_lo = {wire_res_24_65,wire_res_24_64,wire_res_24_63,wire_res_24_62,wire_res_24_61,
    wire_res_24_60,wire_res_24_59,result_reg_r_12_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_12_hi_lo_hi_lo = {wire_res_24_71,wire_res_24_70,wire_res_24_69,wire_res_24_68,wire_res_24_67,
    wire_res_24_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_12_hi_lo = {wire_res_24_78,wire_res_24_77,wire_res_24_76,wire_res_24_75,wire_res_24_74,
    wire_res_24_73,wire_res_24_72,result_reg_r_12_hi_lo_hi_lo,result_reg_r_12_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_12_hi_hi_lo_lo = {wire_res_24_84,wire_res_24_83,wire_res_24_82,wire_res_24_81,wire_res_24_80,
    wire_res_24_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_12_hi_hi_lo = {wire_res_24_91,wire_res_24_90,wire_res_24_89,wire_res_24_88,wire_res_24_87,
    wire_res_24_86,wire_res_24_85,result_reg_r_12_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_12_hi_hi_hi_lo = {wire_res_24_98,wire_res_24_97,wire_res_24_96,wire_res_24_95,wire_res_24_94,
    wire_res_24_93,wire_res_24_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_12_hi = {wire_res_24_105,wire_res_24_104,wire_res_24_103,wire_res_24_102,wire_res_24_101,
    wire_res_24_100,wire_res_24_99,result_reg_r_12_hi_hi_hi_lo,result_reg_r_12_hi_hi_lo,result_reg_r_12_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_12_T = {result_reg_r_12_hi,result_reg_r_12_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [184:0] _a_aux_reg_w_13_T_2 = _GEN_1284 - _T_11288; // @[BinaryDesigns2.scala 225:48]
  wire [184:0] _GEN_52 = wire_res_25_79 ? _a_aux_reg_w_13_T_2 : {{79'd0}, a_aux_reg_r_12}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [183:0] _T_11290 = {b_aux_reg_r_12, 78'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_13 = _GEN_52[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [183:0] _GEN_1363 = {{78'd0}, a_aux_reg_w_13}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_26_78 = _GEN_1363 >= _T_11290; // @[BinaryDesigns2.scala 224:35]
  wire [183:0] _a_aux_reg_r_13_T_2 = _GEN_1363 - _T_11290; // @[BinaryDesigns2.scala 225:48]
  wire [183:0] _GEN_54 = wire_res_26_78 ? _a_aux_reg_r_13_T_2 : {{78'd0}, a_aux_reg_w_13}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_13_lo_lo_lo_lo = {wire_res_26_5,wire_res_26_4,wire_res_26_3,wire_res_26_2,wire_res_26_1,
    wire_res_26_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_13_lo_lo_lo = {wire_res_26_12,wire_res_26_11,wire_res_26_10,wire_res_26_9,wire_res_26_8,
    wire_res_26_7,wire_res_26_6,result_reg_r_13_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_13_lo_lo_hi_lo = {wire_res_26_18,wire_res_26_17,wire_res_26_16,wire_res_26_15,wire_res_26_14,
    wire_res_26_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_13_lo_lo = {wire_res_26_25,wire_res_26_24,wire_res_26_23,wire_res_26_22,wire_res_26_21,
    wire_res_26_20,wire_res_26_19,result_reg_r_13_lo_lo_hi_lo,result_reg_r_13_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_13_lo_hi_lo_lo = {wire_res_26_31,wire_res_26_30,wire_res_26_29,wire_res_26_28,wire_res_26_27,
    wire_res_26_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_13_lo_hi_lo = {wire_res_26_38,wire_res_26_37,wire_res_26_36,wire_res_26_35,wire_res_26_34,
    wire_res_26_33,wire_res_26_32,result_reg_r_13_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_13_lo_hi_hi_lo = {wire_res_26_45,wire_res_26_44,wire_res_26_43,wire_res_26_42,wire_res_26_41,
    wire_res_26_40,wire_res_26_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_13_lo = {wire_res_26_52,wire_res_26_51,wire_res_26_50,wire_res_26_49,wire_res_26_48,
    wire_res_26_47,wire_res_26_46,result_reg_r_13_lo_hi_hi_lo,result_reg_r_13_lo_hi_lo,result_reg_r_13_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_13_hi_lo_lo_lo = {wire_res_26_58,wire_res_26_57,wire_res_26_56,wire_res_26_55,wire_res_26_54,
    wire_res_26_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_13_hi_lo_lo = {wire_res_26_65,wire_res_26_64,wire_res_26_63,wire_res_26_62,wire_res_26_61,
    wire_res_26_60,wire_res_26_59,result_reg_r_13_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_13_hi_lo_hi_lo = {wire_res_26_71,wire_res_26_70,wire_res_26_69,wire_res_26_68,wire_res_26_67,
    wire_res_26_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_13_hi_lo = {wire_res_26_78,wire_res_26_77,wire_res_26_76,wire_res_26_75,wire_res_26_74,
    wire_res_26_73,wire_res_26_72,result_reg_r_13_hi_lo_hi_lo,result_reg_r_13_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_13_hi_hi_lo_lo = {wire_res_26_84,wire_res_26_83,wire_res_26_82,wire_res_26_81,wire_res_26_80,
    wire_res_26_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_13_hi_hi_lo = {wire_res_26_91,wire_res_26_90,wire_res_26_89,wire_res_26_88,wire_res_26_87,
    wire_res_26_86,wire_res_26_85,result_reg_r_13_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_13_hi_hi_hi_lo = {wire_res_26_98,wire_res_26_97,wire_res_26_96,wire_res_26_95,wire_res_26_94,
    wire_res_26_93,wire_res_26_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_13_hi = {wire_res_26_105,wire_res_26_104,wire_res_26_103,wire_res_26_102,wire_res_26_101,
    wire_res_26_100,wire_res_26_99,result_reg_r_13_hi_hi_hi_lo,result_reg_r_13_hi_hi_lo,result_reg_r_13_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_13_T = {result_reg_r_13_hi,result_reg_r_13_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [182:0] _a_aux_reg_w_14_T_2 = _GEN_1285 - _T_11292; // @[BinaryDesigns2.scala 225:48]
  wire [182:0] _GEN_56 = wire_res_27_77 ? _a_aux_reg_w_14_T_2 : {{77'd0}, a_aux_reg_r_13}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [181:0] _T_11294 = {b_aux_reg_r_13, 76'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_14 = _GEN_56[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [181:0] _GEN_1366 = {{76'd0}, a_aux_reg_w_14}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_28_76 = _GEN_1366 >= _T_11294; // @[BinaryDesigns2.scala 224:35]
  wire [181:0] _a_aux_reg_r_14_T_2 = _GEN_1366 - _T_11294; // @[BinaryDesigns2.scala 225:48]
  wire [181:0] _GEN_58 = wire_res_28_76 ? _a_aux_reg_r_14_T_2 : {{76'd0}, a_aux_reg_w_14}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_14_lo_lo_lo_lo = {wire_res_28_5,wire_res_28_4,wire_res_28_3,wire_res_28_2,wire_res_28_1,
    wire_res_28_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_14_lo_lo_lo = {wire_res_28_12,wire_res_28_11,wire_res_28_10,wire_res_28_9,wire_res_28_8,
    wire_res_28_7,wire_res_28_6,result_reg_r_14_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_14_lo_lo_hi_lo = {wire_res_28_18,wire_res_28_17,wire_res_28_16,wire_res_28_15,wire_res_28_14,
    wire_res_28_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_14_lo_lo = {wire_res_28_25,wire_res_28_24,wire_res_28_23,wire_res_28_22,wire_res_28_21,
    wire_res_28_20,wire_res_28_19,result_reg_r_14_lo_lo_hi_lo,result_reg_r_14_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_14_lo_hi_lo_lo = {wire_res_28_31,wire_res_28_30,wire_res_28_29,wire_res_28_28,wire_res_28_27,
    wire_res_28_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_14_lo_hi_lo = {wire_res_28_38,wire_res_28_37,wire_res_28_36,wire_res_28_35,wire_res_28_34,
    wire_res_28_33,wire_res_28_32,result_reg_r_14_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_14_lo_hi_hi_lo = {wire_res_28_45,wire_res_28_44,wire_res_28_43,wire_res_28_42,wire_res_28_41,
    wire_res_28_40,wire_res_28_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_14_lo = {wire_res_28_52,wire_res_28_51,wire_res_28_50,wire_res_28_49,wire_res_28_48,
    wire_res_28_47,wire_res_28_46,result_reg_r_14_lo_hi_hi_lo,result_reg_r_14_lo_hi_lo,result_reg_r_14_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_14_hi_lo_lo_lo = {wire_res_28_58,wire_res_28_57,wire_res_28_56,wire_res_28_55,wire_res_28_54,
    wire_res_28_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_14_hi_lo_lo = {wire_res_28_65,wire_res_28_64,wire_res_28_63,wire_res_28_62,wire_res_28_61,
    wire_res_28_60,wire_res_28_59,result_reg_r_14_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_14_hi_lo_hi_lo = {wire_res_28_71,wire_res_28_70,wire_res_28_69,wire_res_28_68,wire_res_28_67,
    wire_res_28_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_14_hi_lo = {wire_res_28_78,wire_res_28_77,wire_res_28_76,wire_res_28_75,wire_res_28_74,
    wire_res_28_73,wire_res_28_72,result_reg_r_14_hi_lo_hi_lo,result_reg_r_14_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_14_hi_hi_lo_lo = {wire_res_28_84,wire_res_28_83,wire_res_28_82,wire_res_28_81,wire_res_28_80,
    wire_res_28_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_14_hi_hi_lo = {wire_res_28_91,wire_res_28_90,wire_res_28_89,wire_res_28_88,wire_res_28_87,
    wire_res_28_86,wire_res_28_85,result_reg_r_14_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_14_hi_hi_hi_lo = {wire_res_28_98,wire_res_28_97,wire_res_28_96,wire_res_28_95,wire_res_28_94,
    wire_res_28_93,wire_res_28_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_14_hi = {wire_res_28_105,wire_res_28_104,wire_res_28_103,wire_res_28_102,wire_res_28_101,
    wire_res_28_100,wire_res_28_99,result_reg_r_14_hi_hi_hi_lo,result_reg_r_14_hi_hi_lo,result_reg_r_14_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_14_T = {result_reg_r_14_hi,result_reg_r_14_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [180:0] _a_aux_reg_w_15_T_2 = _GEN_1286 - _T_11296; // @[BinaryDesigns2.scala 225:48]
  wire [180:0] _GEN_60 = wire_res_29_75 ? _a_aux_reg_w_15_T_2 : {{75'd0}, a_aux_reg_r_14}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [179:0] _T_11298 = {b_aux_reg_r_14, 74'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_15 = _GEN_60[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [179:0] _GEN_1369 = {{74'd0}, a_aux_reg_w_15}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_30_74 = _GEN_1369 >= _T_11298; // @[BinaryDesigns2.scala 224:35]
  wire [179:0] _a_aux_reg_r_15_T_2 = _GEN_1369 - _T_11298; // @[BinaryDesigns2.scala 225:48]
  wire [179:0] _GEN_62 = wire_res_30_74 ? _a_aux_reg_r_15_T_2 : {{74'd0}, a_aux_reg_w_15}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_15_lo_lo_lo_lo = {wire_res_30_5,wire_res_30_4,wire_res_30_3,wire_res_30_2,wire_res_30_1,
    wire_res_30_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_15_lo_lo_lo = {wire_res_30_12,wire_res_30_11,wire_res_30_10,wire_res_30_9,wire_res_30_8,
    wire_res_30_7,wire_res_30_6,result_reg_r_15_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_15_lo_lo_hi_lo = {wire_res_30_18,wire_res_30_17,wire_res_30_16,wire_res_30_15,wire_res_30_14,
    wire_res_30_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_15_lo_lo = {wire_res_30_25,wire_res_30_24,wire_res_30_23,wire_res_30_22,wire_res_30_21,
    wire_res_30_20,wire_res_30_19,result_reg_r_15_lo_lo_hi_lo,result_reg_r_15_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_15_lo_hi_lo_lo = {wire_res_30_31,wire_res_30_30,wire_res_30_29,wire_res_30_28,wire_res_30_27,
    wire_res_30_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_15_lo_hi_lo = {wire_res_30_38,wire_res_30_37,wire_res_30_36,wire_res_30_35,wire_res_30_34,
    wire_res_30_33,wire_res_30_32,result_reg_r_15_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_15_lo_hi_hi_lo = {wire_res_30_45,wire_res_30_44,wire_res_30_43,wire_res_30_42,wire_res_30_41,
    wire_res_30_40,wire_res_30_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_15_lo = {wire_res_30_52,wire_res_30_51,wire_res_30_50,wire_res_30_49,wire_res_30_48,
    wire_res_30_47,wire_res_30_46,result_reg_r_15_lo_hi_hi_lo,result_reg_r_15_lo_hi_lo,result_reg_r_15_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_15_hi_lo_lo_lo = {wire_res_30_58,wire_res_30_57,wire_res_30_56,wire_res_30_55,wire_res_30_54,
    wire_res_30_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_15_hi_lo_lo = {wire_res_30_65,wire_res_30_64,wire_res_30_63,wire_res_30_62,wire_res_30_61,
    wire_res_30_60,wire_res_30_59,result_reg_r_15_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_15_hi_lo_hi_lo = {wire_res_30_71,wire_res_30_70,wire_res_30_69,wire_res_30_68,wire_res_30_67,
    wire_res_30_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_15_hi_lo = {wire_res_30_78,wire_res_30_77,wire_res_30_76,wire_res_30_75,wire_res_30_74,
    wire_res_30_73,wire_res_30_72,result_reg_r_15_hi_lo_hi_lo,result_reg_r_15_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_15_hi_hi_lo_lo = {wire_res_30_84,wire_res_30_83,wire_res_30_82,wire_res_30_81,wire_res_30_80,
    wire_res_30_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_15_hi_hi_lo = {wire_res_30_91,wire_res_30_90,wire_res_30_89,wire_res_30_88,wire_res_30_87,
    wire_res_30_86,wire_res_30_85,result_reg_r_15_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_15_hi_hi_hi_lo = {wire_res_30_98,wire_res_30_97,wire_res_30_96,wire_res_30_95,wire_res_30_94,
    wire_res_30_93,wire_res_30_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_15_hi = {wire_res_30_105,wire_res_30_104,wire_res_30_103,wire_res_30_102,wire_res_30_101,
    wire_res_30_100,wire_res_30_99,result_reg_r_15_hi_hi_hi_lo,result_reg_r_15_hi_hi_lo,result_reg_r_15_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_15_T = {result_reg_r_15_hi,result_reg_r_15_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [178:0] _a_aux_reg_w_16_T_2 = _GEN_1287 - _T_11300; // @[BinaryDesigns2.scala 225:48]
  wire [178:0] _GEN_64 = wire_res_31_73 ? _a_aux_reg_w_16_T_2 : {{73'd0}, a_aux_reg_r_15}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [177:0] _T_11302 = {b_aux_reg_r_15, 72'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_16 = _GEN_64[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [177:0] _GEN_1372 = {{72'd0}, a_aux_reg_w_16}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_32_72 = _GEN_1372 >= _T_11302; // @[BinaryDesigns2.scala 224:35]
  wire [177:0] _a_aux_reg_r_16_T_2 = _GEN_1372 - _T_11302; // @[BinaryDesigns2.scala 225:48]
  wire [177:0] _GEN_66 = wire_res_32_72 ? _a_aux_reg_r_16_T_2 : {{72'd0}, a_aux_reg_w_16}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_16_lo_lo_lo_lo = {wire_res_32_5,wire_res_32_4,wire_res_32_3,wire_res_32_2,wire_res_32_1,
    wire_res_32_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_16_lo_lo_lo = {wire_res_32_12,wire_res_32_11,wire_res_32_10,wire_res_32_9,wire_res_32_8,
    wire_res_32_7,wire_res_32_6,result_reg_r_16_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_16_lo_lo_hi_lo = {wire_res_32_18,wire_res_32_17,wire_res_32_16,wire_res_32_15,wire_res_32_14,
    wire_res_32_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_16_lo_lo = {wire_res_32_25,wire_res_32_24,wire_res_32_23,wire_res_32_22,wire_res_32_21,
    wire_res_32_20,wire_res_32_19,result_reg_r_16_lo_lo_hi_lo,result_reg_r_16_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_16_lo_hi_lo_lo = {wire_res_32_31,wire_res_32_30,wire_res_32_29,wire_res_32_28,wire_res_32_27,
    wire_res_32_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_16_lo_hi_lo = {wire_res_32_38,wire_res_32_37,wire_res_32_36,wire_res_32_35,wire_res_32_34,
    wire_res_32_33,wire_res_32_32,result_reg_r_16_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_16_lo_hi_hi_lo = {wire_res_32_45,wire_res_32_44,wire_res_32_43,wire_res_32_42,wire_res_32_41,
    wire_res_32_40,wire_res_32_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_16_lo = {wire_res_32_52,wire_res_32_51,wire_res_32_50,wire_res_32_49,wire_res_32_48,
    wire_res_32_47,wire_res_32_46,result_reg_r_16_lo_hi_hi_lo,result_reg_r_16_lo_hi_lo,result_reg_r_16_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_16_hi_lo_lo_lo = {wire_res_32_58,wire_res_32_57,wire_res_32_56,wire_res_32_55,wire_res_32_54,
    wire_res_32_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_16_hi_lo_lo = {wire_res_32_65,wire_res_32_64,wire_res_32_63,wire_res_32_62,wire_res_32_61,
    wire_res_32_60,wire_res_32_59,result_reg_r_16_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_16_hi_lo_hi_lo = {wire_res_32_71,wire_res_32_70,wire_res_32_69,wire_res_32_68,wire_res_32_67,
    wire_res_32_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_16_hi_lo = {wire_res_32_78,wire_res_32_77,wire_res_32_76,wire_res_32_75,wire_res_32_74,
    wire_res_32_73,wire_res_32_72,result_reg_r_16_hi_lo_hi_lo,result_reg_r_16_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_16_hi_hi_lo_lo = {wire_res_32_84,wire_res_32_83,wire_res_32_82,wire_res_32_81,wire_res_32_80,
    wire_res_32_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_16_hi_hi_lo = {wire_res_32_91,wire_res_32_90,wire_res_32_89,wire_res_32_88,wire_res_32_87,
    wire_res_32_86,wire_res_32_85,result_reg_r_16_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_16_hi_hi_hi_lo = {wire_res_32_98,wire_res_32_97,wire_res_32_96,wire_res_32_95,wire_res_32_94,
    wire_res_32_93,wire_res_32_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_16_hi = {wire_res_32_105,wire_res_32_104,wire_res_32_103,wire_res_32_102,wire_res_32_101,
    wire_res_32_100,wire_res_32_99,result_reg_r_16_hi_hi_hi_lo,result_reg_r_16_hi_hi_lo,result_reg_r_16_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_16_T = {result_reg_r_16_hi,result_reg_r_16_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [176:0] _a_aux_reg_w_17_T_2 = _GEN_1288 - _T_11304; // @[BinaryDesigns2.scala 225:48]
  wire [176:0] _GEN_68 = wire_res_33_71 ? _a_aux_reg_w_17_T_2 : {{71'd0}, a_aux_reg_r_16}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [175:0] _T_11306 = {b_aux_reg_r_16, 70'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_17 = _GEN_68[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [175:0] _GEN_1375 = {{70'd0}, a_aux_reg_w_17}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_34_70 = _GEN_1375 >= _T_11306; // @[BinaryDesigns2.scala 224:35]
  wire [175:0] _a_aux_reg_r_17_T_2 = _GEN_1375 - _T_11306; // @[BinaryDesigns2.scala 225:48]
  wire [175:0] _GEN_70 = wire_res_34_70 ? _a_aux_reg_r_17_T_2 : {{70'd0}, a_aux_reg_w_17}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_17_lo_lo_lo_lo = {wire_res_34_5,wire_res_34_4,wire_res_34_3,wire_res_34_2,wire_res_34_1,
    wire_res_34_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_17_lo_lo_lo = {wire_res_34_12,wire_res_34_11,wire_res_34_10,wire_res_34_9,wire_res_34_8,
    wire_res_34_7,wire_res_34_6,result_reg_r_17_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_17_lo_lo_hi_lo = {wire_res_34_18,wire_res_34_17,wire_res_34_16,wire_res_34_15,wire_res_34_14,
    wire_res_34_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_17_lo_lo = {wire_res_34_25,wire_res_34_24,wire_res_34_23,wire_res_34_22,wire_res_34_21,
    wire_res_34_20,wire_res_34_19,result_reg_r_17_lo_lo_hi_lo,result_reg_r_17_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_17_lo_hi_lo_lo = {wire_res_34_31,wire_res_34_30,wire_res_34_29,wire_res_34_28,wire_res_34_27,
    wire_res_34_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_17_lo_hi_lo = {wire_res_34_38,wire_res_34_37,wire_res_34_36,wire_res_34_35,wire_res_34_34,
    wire_res_34_33,wire_res_34_32,result_reg_r_17_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_17_lo_hi_hi_lo = {wire_res_34_45,wire_res_34_44,wire_res_34_43,wire_res_34_42,wire_res_34_41,
    wire_res_34_40,wire_res_34_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_17_lo = {wire_res_34_52,wire_res_34_51,wire_res_34_50,wire_res_34_49,wire_res_34_48,
    wire_res_34_47,wire_res_34_46,result_reg_r_17_lo_hi_hi_lo,result_reg_r_17_lo_hi_lo,result_reg_r_17_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_17_hi_lo_lo_lo = {wire_res_34_58,wire_res_34_57,wire_res_34_56,wire_res_34_55,wire_res_34_54,
    wire_res_34_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_17_hi_lo_lo = {wire_res_34_65,wire_res_34_64,wire_res_34_63,wire_res_34_62,wire_res_34_61,
    wire_res_34_60,wire_res_34_59,result_reg_r_17_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_17_hi_lo_hi_lo = {wire_res_34_71,wire_res_34_70,wire_res_34_69,wire_res_34_68,wire_res_34_67,
    wire_res_34_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_17_hi_lo = {wire_res_34_78,wire_res_34_77,wire_res_34_76,wire_res_34_75,wire_res_34_74,
    wire_res_34_73,wire_res_34_72,result_reg_r_17_hi_lo_hi_lo,result_reg_r_17_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_17_hi_hi_lo_lo = {wire_res_34_84,wire_res_34_83,wire_res_34_82,wire_res_34_81,wire_res_34_80,
    wire_res_34_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_17_hi_hi_lo = {wire_res_34_91,wire_res_34_90,wire_res_34_89,wire_res_34_88,wire_res_34_87,
    wire_res_34_86,wire_res_34_85,result_reg_r_17_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_17_hi_hi_hi_lo = {wire_res_34_98,wire_res_34_97,wire_res_34_96,wire_res_34_95,wire_res_34_94,
    wire_res_34_93,wire_res_34_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_17_hi = {wire_res_34_105,wire_res_34_104,wire_res_34_103,wire_res_34_102,wire_res_34_101,
    wire_res_34_100,wire_res_34_99,result_reg_r_17_hi_hi_hi_lo,result_reg_r_17_hi_hi_lo,result_reg_r_17_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_17_T = {result_reg_r_17_hi,result_reg_r_17_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [174:0] _a_aux_reg_w_18_T_2 = _GEN_1289 - _T_11308; // @[BinaryDesigns2.scala 225:48]
  wire [174:0] _GEN_72 = wire_res_35_69 ? _a_aux_reg_w_18_T_2 : {{69'd0}, a_aux_reg_r_17}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [173:0] _T_11310 = {b_aux_reg_r_17, 68'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_18 = _GEN_72[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [173:0] _GEN_1378 = {{68'd0}, a_aux_reg_w_18}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_36_68 = _GEN_1378 >= _T_11310; // @[BinaryDesigns2.scala 224:35]
  wire [173:0] _a_aux_reg_r_18_T_2 = _GEN_1378 - _T_11310; // @[BinaryDesigns2.scala 225:48]
  wire [173:0] _GEN_74 = wire_res_36_68 ? _a_aux_reg_r_18_T_2 : {{68'd0}, a_aux_reg_w_18}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_18_lo_lo_lo_lo = {wire_res_36_5,wire_res_36_4,wire_res_36_3,wire_res_36_2,wire_res_36_1,
    wire_res_36_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_18_lo_lo_lo = {wire_res_36_12,wire_res_36_11,wire_res_36_10,wire_res_36_9,wire_res_36_8,
    wire_res_36_7,wire_res_36_6,result_reg_r_18_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_18_lo_lo_hi_lo = {wire_res_36_18,wire_res_36_17,wire_res_36_16,wire_res_36_15,wire_res_36_14,
    wire_res_36_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_18_lo_lo = {wire_res_36_25,wire_res_36_24,wire_res_36_23,wire_res_36_22,wire_res_36_21,
    wire_res_36_20,wire_res_36_19,result_reg_r_18_lo_lo_hi_lo,result_reg_r_18_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_18_lo_hi_lo_lo = {wire_res_36_31,wire_res_36_30,wire_res_36_29,wire_res_36_28,wire_res_36_27,
    wire_res_36_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_18_lo_hi_lo = {wire_res_36_38,wire_res_36_37,wire_res_36_36,wire_res_36_35,wire_res_36_34,
    wire_res_36_33,wire_res_36_32,result_reg_r_18_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_18_lo_hi_hi_lo = {wire_res_36_45,wire_res_36_44,wire_res_36_43,wire_res_36_42,wire_res_36_41,
    wire_res_36_40,wire_res_36_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_18_lo = {wire_res_36_52,wire_res_36_51,wire_res_36_50,wire_res_36_49,wire_res_36_48,
    wire_res_36_47,wire_res_36_46,result_reg_r_18_lo_hi_hi_lo,result_reg_r_18_lo_hi_lo,result_reg_r_18_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_18_hi_lo_lo_lo = {wire_res_36_58,wire_res_36_57,wire_res_36_56,wire_res_36_55,wire_res_36_54,
    wire_res_36_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_18_hi_lo_lo = {wire_res_36_65,wire_res_36_64,wire_res_36_63,wire_res_36_62,wire_res_36_61,
    wire_res_36_60,wire_res_36_59,result_reg_r_18_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_18_hi_lo_hi_lo = {wire_res_36_71,wire_res_36_70,wire_res_36_69,wire_res_36_68,wire_res_36_67,
    wire_res_36_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_18_hi_lo = {wire_res_36_78,wire_res_36_77,wire_res_36_76,wire_res_36_75,wire_res_36_74,
    wire_res_36_73,wire_res_36_72,result_reg_r_18_hi_lo_hi_lo,result_reg_r_18_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_18_hi_hi_lo_lo = {wire_res_36_84,wire_res_36_83,wire_res_36_82,wire_res_36_81,wire_res_36_80,
    wire_res_36_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_18_hi_hi_lo = {wire_res_36_91,wire_res_36_90,wire_res_36_89,wire_res_36_88,wire_res_36_87,
    wire_res_36_86,wire_res_36_85,result_reg_r_18_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_18_hi_hi_hi_lo = {wire_res_36_98,wire_res_36_97,wire_res_36_96,wire_res_36_95,wire_res_36_94,
    wire_res_36_93,wire_res_36_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_18_hi = {wire_res_36_105,wire_res_36_104,wire_res_36_103,wire_res_36_102,wire_res_36_101,
    wire_res_36_100,wire_res_36_99,result_reg_r_18_hi_hi_hi_lo,result_reg_r_18_hi_hi_lo,result_reg_r_18_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_18_T = {result_reg_r_18_hi,result_reg_r_18_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [172:0] _a_aux_reg_w_19_T_2 = _GEN_1290 - _T_11312; // @[BinaryDesigns2.scala 225:48]
  wire [172:0] _GEN_76 = wire_res_37_67 ? _a_aux_reg_w_19_T_2 : {{67'd0}, a_aux_reg_r_18}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [171:0] _T_11314 = {b_aux_reg_r_18, 66'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_19 = _GEN_76[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [171:0] _GEN_1381 = {{66'd0}, a_aux_reg_w_19}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_38_66 = _GEN_1381 >= _T_11314; // @[BinaryDesigns2.scala 224:35]
  wire [171:0] _a_aux_reg_r_19_T_2 = _GEN_1381 - _T_11314; // @[BinaryDesigns2.scala 225:48]
  wire [171:0] _GEN_78 = wire_res_38_66 ? _a_aux_reg_r_19_T_2 : {{66'd0}, a_aux_reg_w_19}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_19_lo_lo_lo_lo = {wire_res_38_5,wire_res_38_4,wire_res_38_3,wire_res_38_2,wire_res_38_1,
    wire_res_38_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_19_lo_lo_lo = {wire_res_38_12,wire_res_38_11,wire_res_38_10,wire_res_38_9,wire_res_38_8,
    wire_res_38_7,wire_res_38_6,result_reg_r_19_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_19_lo_lo_hi_lo = {wire_res_38_18,wire_res_38_17,wire_res_38_16,wire_res_38_15,wire_res_38_14,
    wire_res_38_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_19_lo_lo = {wire_res_38_25,wire_res_38_24,wire_res_38_23,wire_res_38_22,wire_res_38_21,
    wire_res_38_20,wire_res_38_19,result_reg_r_19_lo_lo_hi_lo,result_reg_r_19_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_19_lo_hi_lo_lo = {wire_res_38_31,wire_res_38_30,wire_res_38_29,wire_res_38_28,wire_res_38_27,
    wire_res_38_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_19_lo_hi_lo = {wire_res_38_38,wire_res_38_37,wire_res_38_36,wire_res_38_35,wire_res_38_34,
    wire_res_38_33,wire_res_38_32,result_reg_r_19_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_19_lo_hi_hi_lo = {wire_res_38_45,wire_res_38_44,wire_res_38_43,wire_res_38_42,wire_res_38_41,
    wire_res_38_40,wire_res_38_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_19_lo = {wire_res_38_52,wire_res_38_51,wire_res_38_50,wire_res_38_49,wire_res_38_48,
    wire_res_38_47,wire_res_38_46,result_reg_r_19_lo_hi_hi_lo,result_reg_r_19_lo_hi_lo,result_reg_r_19_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_19_hi_lo_lo_lo = {wire_res_38_58,wire_res_38_57,wire_res_38_56,wire_res_38_55,wire_res_38_54,
    wire_res_38_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_19_hi_lo_lo = {wire_res_38_65,wire_res_38_64,wire_res_38_63,wire_res_38_62,wire_res_38_61,
    wire_res_38_60,wire_res_38_59,result_reg_r_19_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_19_hi_lo_hi_lo = {wire_res_38_71,wire_res_38_70,wire_res_38_69,wire_res_38_68,wire_res_38_67,
    wire_res_38_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_19_hi_lo = {wire_res_38_78,wire_res_38_77,wire_res_38_76,wire_res_38_75,wire_res_38_74,
    wire_res_38_73,wire_res_38_72,result_reg_r_19_hi_lo_hi_lo,result_reg_r_19_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_19_hi_hi_lo_lo = {wire_res_38_84,wire_res_38_83,wire_res_38_82,wire_res_38_81,wire_res_38_80,
    wire_res_38_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_19_hi_hi_lo = {wire_res_38_91,wire_res_38_90,wire_res_38_89,wire_res_38_88,wire_res_38_87,
    wire_res_38_86,wire_res_38_85,result_reg_r_19_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_19_hi_hi_hi_lo = {wire_res_38_98,wire_res_38_97,wire_res_38_96,wire_res_38_95,wire_res_38_94,
    wire_res_38_93,wire_res_38_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_19_hi = {wire_res_38_105,wire_res_38_104,wire_res_38_103,wire_res_38_102,wire_res_38_101,
    wire_res_38_100,wire_res_38_99,result_reg_r_19_hi_hi_hi_lo,result_reg_r_19_hi_hi_lo,result_reg_r_19_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_19_T = {result_reg_r_19_hi,result_reg_r_19_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [170:0] _a_aux_reg_w_20_T_2 = _GEN_1291 - _T_11316; // @[BinaryDesigns2.scala 225:48]
  wire [170:0] _GEN_80 = wire_res_39_65 ? _a_aux_reg_w_20_T_2 : {{65'd0}, a_aux_reg_r_19}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [169:0] _T_11318 = {b_aux_reg_r_19, 64'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_20 = _GEN_80[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [169:0] _GEN_1384 = {{64'd0}, a_aux_reg_w_20}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_40_64 = _GEN_1384 >= _T_11318; // @[BinaryDesigns2.scala 224:35]
  wire [169:0] _a_aux_reg_r_20_T_2 = _GEN_1384 - _T_11318; // @[BinaryDesigns2.scala 225:48]
  wire [169:0] _GEN_82 = wire_res_40_64 ? _a_aux_reg_r_20_T_2 : {{64'd0}, a_aux_reg_w_20}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_20_lo_lo_lo_lo = {wire_res_40_5,wire_res_40_4,wire_res_40_3,wire_res_40_2,wire_res_40_1,
    wire_res_40_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_20_lo_lo_lo = {wire_res_40_12,wire_res_40_11,wire_res_40_10,wire_res_40_9,wire_res_40_8,
    wire_res_40_7,wire_res_40_6,result_reg_r_20_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_20_lo_lo_hi_lo = {wire_res_40_18,wire_res_40_17,wire_res_40_16,wire_res_40_15,wire_res_40_14,
    wire_res_40_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_20_lo_lo = {wire_res_40_25,wire_res_40_24,wire_res_40_23,wire_res_40_22,wire_res_40_21,
    wire_res_40_20,wire_res_40_19,result_reg_r_20_lo_lo_hi_lo,result_reg_r_20_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_20_lo_hi_lo_lo = {wire_res_40_31,wire_res_40_30,wire_res_40_29,wire_res_40_28,wire_res_40_27,
    wire_res_40_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_20_lo_hi_lo = {wire_res_40_38,wire_res_40_37,wire_res_40_36,wire_res_40_35,wire_res_40_34,
    wire_res_40_33,wire_res_40_32,result_reg_r_20_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_20_lo_hi_hi_lo = {wire_res_40_45,wire_res_40_44,wire_res_40_43,wire_res_40_42,wire_res_40_41,
    wire_res_40_40,wire_res_40_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_20_lo = {wire_res_40_52,wire_res_40_51,wire_res_40_50,wire_res_40_49,wire_res_40_48,
    wire_res_40_47,wire_res_40_46,result_reg_r_20_lo_hi_hi_lo,result_reg_r_20_lo_hi_lo,result_reg_r_20_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_20_hi_lo_lo_lo = {wire_res_40_58,wire_res_40_57,wire_res_40_56,wire_res_40_55,wire_res_40_54,
    wire_res_40_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_20_hi_lo_lo = {wire_res_40_65,wire_res_40_64,wire_res_40_63,wire_res_40_62,wire_res_40_61,
    wire_res_40_60,wire_res_40_59,result_reg_r_20_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_20_hi_lo_hi_lo = {wire_res_40_71,wire_res_40_70,wire_res_40_69,wire_res_40_68,wire_res_40_67,
    wire_res_40_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_20_hi_lo = {wire_res_40_78,wire_res_40_77,wire_res_40_76,wire_res_40_75,wire_res_40_74,
    wire_res_40_73,wire_res_40_72,result_reg_r_20_hi_lo_hi_lo,result_reg_r_20_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_20_hi_hi_lo_lo = {wire_res_40_84,wire_res_40_83,wire_res_40_82,wire_res_40_81,wire_res_40_80,
    wire_res_40_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_20_hi_hi_lo = {wire_res_40_91,wire_res_40_90,wire_res_40_89,wire_res_40_88,wire_res_40_87,
    wire_res_40_86,wire_res_40_85,result_reg_r_20_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_20_hi_hi_hi_lo = {wire_res_40_98,wire_res_40_97,wire_res_40_96,wire_res_40_95,wire_res_40_94,
    wire_res_40_93,wire_res_40_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_20_hi = {wire_res_40_105,wire_res_40_104,wire_res_40_103,wire_res_40_102,wire_res_40_101,
    wire_res_40_100,wire_res_40_99,result_reg_r_20_hi_hi_hi_lo,result_reg_r_20_hi_hi_lo,result_reg_r_20_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_20_T = {result_reg_r_20_hi,result_reg_r_20_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [168:0] _a_aux_reg_w_21_T_2 = _GEN_1292 - _T_11320; // @[BinaryDesigns2.scala 225:48]
  wire [168:0] _GEN_84 = wire_res_41_63 ? _a_aux_reg_w_21_T_2 : {{63'd0}, a_aux_reg_r_20}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [167:0] _T_11322 = {b_aux_reg_r_20, 62'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_21 = _GEN_84[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [167:0] _GEN_1387 = {{62'd0}, a_aux_reg_w_21}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_42_62 = _GEN_1387 >= _T_11322; // @[BinaryDesigns2.scala 224:35]
  wire [167:0] _a_aux_reg_r_21_T_2 = _GEN_1387 - _T_11322; // @[BinaryDesigns2.scala 225:48]
  wire [167:0] _GEN_86 = wire_res_42_62 ? _a_aux_reg_r_21_T_2 : {{62'd0}, a_aux_reg_w_21}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_21_lo_lo_lo_lo = {wire_res_42_5,wire_res_42_4,wire_res_42_3,wire_res_42_2,wire_res_42_1,
    wire_res_42_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_21_lo_lo_lo = {wire_res_42_12,wire_res_42_11,wire_res_42_10,wire_res_42_9,wire_res_42_8,
    wire_res_42_7,wire_res_42_6,result_reg_r_21_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_21_lo_lo_hi_lo = {wire_res_42_18,wire_res_42_17,wire_res_42_16,wire_res_42_15,wire_res_42_14,
    wire_res_42_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_21_lo_lo = {wire_res_42_25,wire_res_42_24,wire_res_42_23,wire_res_42_22,wire_res_42_21,
    wire_res_42_20,wire_res_42_19,result_reg_r_21_lo_lo_hi_lo,result_reg_r_21_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_21_lo_hi_lo_lo = {wire_res_42_31,wire_res_42_30,wire_res_42_29,wire_res_42_28,wire_res_42_27,
    wire_res_42_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_21_lo_hi_lo = {wire_res_42_38,wire_res_42_37,wire_res_42_36,wire_res_42_35,wire_res_42_34,
    wire_res_42_33,wire_res_42_32,result_reg_r_21_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_21_lo_hi_hi_lo = {wire_res_42_45,wire_res_42_44,wire_res_42_43,wire_res_42_42,wire_res_42_41,
    wire_res_42_40,wire_res_42_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_21_lo = {wire_res_42_52,wire_res_42_51,wire_res_42_50,wire_res_42_49,wire_res_42_48,
    wire_res_42_47,wire_res_42_46,result_reg_r_21_lo_hi_hi_lo,result_reg_r_21_lo_hi_lo,result_reg_r_21_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_21_hi_lo_lo_lo = {wire_res_42_58,wire_res_42_57,wire_res_42_56,wire_res_42_55,wire_res_42_54,
    wire_res_42_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_21_hi_lo_lo = {wire_res_42_65,wire_res_42_64,wire_res_42_63,wire_res_42_62,wire_res_42_61,
    wire_res_42_60,wire_res_42_59,result_reg_r_21_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_21_hi_lo_hi_lo = {wire_res_42_71,wire_res_42_70,wire_res_42_69,wire_res_42_68,wire_res_42_67,
    wire_res_42_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_21_hi_lo = {wire_res_42_78,wire_res_42_77,wire_res_42_76,wire_res_42_75,wire_res_42_74,
    wire_res_42_73,wire_res_42_72,result_reg_r_21_hi_lo_hi_lo,result_reg_r_21_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_21_hi_hi_lo_lo = {wire_res_42_84,wire_res_42_83,wire_res_42_82,wire_res_42_81,wire_res_42_80,
    wire_res_42_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_21_hi_hi_lo = {wire_res_42_91,wire_res_42_90,wire_res_42_89,wire_res_42_88,wire_res_42_87,
    wire_res_42_86,wire_res_42_85,result_reg_r_21_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_21_hi_hi_hi_lo = {wire_res_42_98,wire_res_42_97,wire_res_42_96,wire_res_42_95,wire_res_42_94,
    wire_res_42_93,wire_res_42_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_21_hi = {wire_res_42_105,wire_res_42_104,wire_res_42_103,wire_res_42_102,wire_res_42_101,
    wire_res_42_100,wire_res_42_99,result_reg_r_21_hi_hi_hi_lo,result_reg_r_21_hi_hi_lo,result_reg_r_21_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_21_T = {result_reg_r_21_hi,result_reg_r_21_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [166:0] _a_aux_reg_w_22_T_2 = _GEN_1293 - _T_11324; // @[BinaryDesigns2.scala 225:48]
  wire [166:0] _GEN_88 = wire_res_43_61 ? _a_aux_reg_w_22_T_2 : {{61'd0}, a_aux_reg_r_21}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [165:0] _T_11326 = {b_aux_reg_r_21, 60'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_22 = _GEN_88[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [165:0] _GEN_1390 = {{60'd0}, a_aux_reg_w_22}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_44_60 = _GEN_1390 >= _T_11326; // @[BinaryDesigns2.scala 224:35]
  wire [165:0] _a_aux_reg_r_22_T_2 = _GEN_1390 - _T_11326; // @[BinaryDesigns2.scala 225:48]
  wire [165:0] _GEN_90 = wire_res_44_60 ? _a_aux_reg_r_22_T_2 : {{60'd0}, a_aux_reg_w_22}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_22_lo_lo_lo_lo = {wire_res_44_5,wire_res_44_4,wire_res_44_3,wire_res_44_2,wire_res_44_1,
    wire_res_44_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_22_lo_lo_lo = {wire_res_44_12,wire_res_44_11,wire_res_44_10,wire_res_44_9,wire_res_44_8,
    wire_res_44_7,wire_res_44_6,result_reg_r_22_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_22_lo_lo_hi_lo = {wire_res_44_18,wire_res_44_17,wire_res_44_16,wire_res_44_15,wire_res_44_14,
    wire_res_44_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_22_lo_lo = {wire_res_44_25,wire_res_44_24,wire_res_44_23,wire_res_44_22,wire_res_44_21,
    wire_res_44_20,wire_res_44_19,result_reg_r_22_lo_lo_hi_lo,result_reg_r_22_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_22_lo_hi_lo_lo = {wire_res_44_31,wire_res_44_30,wire_res_44_29,wire_res_44_28,wire_res_44_27,
    wire_res_44_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_22_lo_hi_lo = {wire_res_44_38,wire_res_44_37,wire_res_44_36,wire_res_44_35,wire_res_44_34,
    wire_res_44_33,wire_res_44_32,result_reg_r_22_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_22_lo_hi_hi_lo = {wire_res_44_45,wire_res_44_44,wire_res_44_43,wire_res_44_42,wire_res_44_41,
    wire_res_44_40,wire_res_44_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_22_lo = {wire_res_44_52,wire_res_44_51,wire_res_44_50,wire_res_44_49,wire_res_44_48,
    wire_res_44_47,wire_res_44_46,result_reg_r_22_lo_hi_hi_lo,result_reg_r_22_lo_hi_lo,result_reg_r_22_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_22_hi_lo_lo_lo = {wire_res_44_58,wire_res_44_57,wire_res_44_56,wire_res_44_55,wire_res_44_54,
    wire_res_44_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_22_hi_lo_lo = {wire_res_44_65,wire_res_44_64,wire_res_44_63,wire_res_44_62,wire_res_44_61,
    wire_res_44_60,wire_res_44_59,result_reg_r_22_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_22_hi_lo_hi_lo = {wire_res_44_71,wire_res_44_70,wire_res_44_69,wire_res_44_68,wire_res_44_67,
    wire_res_44_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_22_hi_lo = {wire_res_44_78,wire_res_44_77,wire_res_44_76,wire_res_44_75,wire_res_44_74,
    wire_res_44_73,wire_res_44_72,result_reg_r_22_hi_lo_hi_lo,result_reg_r_22_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_22_hi_hi_lo_lo = {wire_res_44_84,wire_res_44_83,wire_res_44_82,wire_res_44_81,wire_res_44_80,
    wire_res_44_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_22_hi_hi_lo = {wire_res_44_91,wire_res_44_90,wire_res_44_89,wire_res_44_88,wire_res_44_87,
    wire_res_44_86,wire_res_44_85,result_reg_r_22_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_22_hi_hi_hi_lo = {wire_res_44_98,wire_res_44_97,wire_res_44_96,wire_res_44_95,wire_res_44_94,
    wire_res_44_93,wire_res_44_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_22_hi = {wire_res_44_105,wire_res_44_104,wire_res_44_103,wire_res_44_102,wire_res_44_101,
    wire_res_44_100,wire_res_44_99,result_reg_r_22_hi_hi_hi_lo,result_reg_r_22_hi_hi_lo,result_reg_r_22_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_22_T = {result_reg_r_22_hi,result_reg_r_22_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [164:0] _a_aux_reg_w_23_T_2 = _GEN_1294 - _T_11328; // @[BinaryDesigns2.scala 225:48]
  wire [164:0] _GEN_92 = wire_res_45_59 ? _a_aux_reg_w_23_T_2 : {{59'd0}, a_aux_reg_r_22}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [163:0] _T_11330 = {b_aux_reg_r_22, 58'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_23 = _GEN_92[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [163:0] _GEN_1393 = {{58'd0}, a_aux_reg_w_23}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_46_58 = _GEN_1393 >= _T_11330; // @[BinaryDesigns2.scala 224:35]
  wire [163:0] _a_aux_reg_r_23_T_2 = _GEN_1393 - _T_11330; // @[BinaryDesigns2.scala 225:48]
  wire [163:0] _GEN_94 = wire_res_46_58 ? _a_aux_reg_r_23_T_2 : {{58'd0}, a_aux_reg_w_23}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_23_lo_lo_lo_lo = {wire_res_46_5,wire_res_46_4,wire_res_46_3,wire_res_46_2,wire_res_46_1,
    wire_res_46_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_23_lo_lo_lo = {wire_res_46_12,wire_res_46_11,wire_res_46_10,wire_res_46_9,wire_res_46_8,
    wire_res_46_7,wire_res_46_6,result_reg_r_23_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_23_lo_lo_hi_lo = {wire_res_46_18,wire_res_46_17,wire_res_46_16,wire_res_46_15,wire_res_46_14,
    wire_res_46_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_23_lo_lo = {wire_res_46_25,wire_res_46_24,wire_res_46_23,wire_res_46_22,wire_res_46_21,
    wire_res_46_20,wire_res_46_19,result_reg_r_23_lo_lo_hi_lo,result_reg_r_23_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_23_lo_hi_lo_lo = {wire_res_46_31,wire_res_46_30,wire_res_46_29,wire_res_46_28,wire_res_46_27,
    wire_res_46_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_23_lo_hi_lo = {wire_res_46_38,wire_res_46_37,wire_res_46_36,wire_res_46_35,wire_res_46_34,
    wire_res_46_33,wire_res_46_32,result_reg_r_23_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_23_lo_hi_hi_lo = {wire_res_46_45,wire_res_46_44,wire_res_46_43,wire_res_46_42,wire_res_46_41,
    wire_res_46_40,wire_res_46_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_23_lo = {wire_res_46_52,wire_res_46_51,wire_res_46_50,wire_res_46_49,wire_res_46_48,
    wire_res_46_47,wire_res_46_46,result_reg_r_23_lo_hi_hi_lo,result_reg_r_23_lo_hi_lo,result_reg_r_23_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_23_hi_lo_lo_lo = {wire_res_46_58,wire_res_46_57,wire_res_46_56,wire_res_46_55,wire_res_46_54,
    wire_res_46_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_23_hi_lo_lo = {wire_res_46_65,wire_res_46_64,wire_res_46_63,wire_res_46_62,wire_res_46_61,
    wire_res_46_60,wire_res_46_59,result_reg_r_23_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_23_hi_lo_hi_lo = {wire_res_46_71,wire_res_46_70,wire_res_46_69,wire_res_46_68,wire_res_46_67,
    wire_res_46_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_23_hi_lo = {wire_res_46_78,wire_res_46_77,wire_res_46_76,wire_res_46_75,wire_res_46_74,
    wire_res_46_73,wire_res_46_72,result_reg_r_23_hi_lo_hi_lo,result_reg_r_23_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_23_hi_hi_lo_lo = {wire_res_46_84,wire_res_46_83,wire_res_46_82,wire_res_46_81,wire_res_46_80,
    wire_res_46_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_23_hi_hi_lo = {wire_res_46_91,wire_res_46_90,wire_res_46_89,wire_res_46_88,wire_res_46_87,
    wire_res_46_86,wire_res_46_85,result_reg_r_23_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_23_hi_hi_hi_lo = {wire_res_46_98,wire_res_46_97,wire_res_46_96,wire_res_46_95,wire_res_46_94,
    wire_res_46_93,wire_res_46_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_23_hi = {wire_res_46_105,wire_res_46_104,wire_res_46_103,wire_res_46_102,wire_res_46_101,
    wire_res_46_100,wire_res_46_99,result_reg_r_23_hi_hi_hi_lo,result_reg_r_23_hi_hi_lo,result_reg_r_23_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_23_T = {result_reg_r_23_hi,result_reg_r_23_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [162:0] _a_aux_reg_w_24_T_2 = _GEN_1295 - _T_11332; // @[BinaryDesigns2.scala 225:48]
  wire [162:0] _GEN_96 = wire_res_47_57 ? _a_aux_reg_w_24_T_2 : {{57'd0}, a_aux_reg_r_23}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [161:0] _T_11334 = {b_aux_reg_r_23, 56'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_24 = _GEN_96[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [161:0] _GEN_1396 = {{56'd0}, a_aux_reg_w_24}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_48_56 = _GEN_1396 >= _T_11334; // @[BinaryDesigns2.scala 224:35]
  wire [161:0] _a_aux_reg_r_24_T_2 = _GEN_1396 - _T_11334; // @[BinaryDesigns2.scala 225:48]
  wire [161:0] _GEN_98 = wire_res_48_56 ? _a_aux_reg_r_24_T_2 : {{56'd0}, a_aux_reg_w_24}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_24_lo_lo_lo_lo = {wire_res_48_5,wire_res_48_4,wire_res_48_3,wire_res_48_2,wire_res_48_1,
    wire_res_48_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_24_lo_lo_lo = {wire_res_48_12,wire_res_48_11,wire_res_48_10,wire_res_48_9,wire_res_48_8,
    wire_res_48_7,wire_res_48_6,result_reg_r_24_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_24_lo_lo_hi_lo = {wire_res_48_18,wire_res_48_17,wire_res_48_16,wire_res_48_15,wire_res_48_14,
    wire_res_48_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_24_lo_lo = {wire_res_48_25,wire_res_48_24,wire_res_48_23,wire_res_48_22,wire_res_48_21,
    wire_res_48_20,wire_res_48_19,result_reg_r_24_lo_lo_hi_lo,result_reg_r_24_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_24_lo_hi_lo_lo = {wire_res_48_31,wire_res_48_30,wire_res_48_29,wire_res_48_28,wire_res_48_27,
    wire_res_48_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_24_lo_hi_lo = {wire_res_48_38,wire_res_48_37,wire_res_48_36,wire_res_48_35,wire_res_48_34,
    wire_res_48_33,wire_res_48_32,result_reg_r_24_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_24_lo_hi_hi_lo = {wire_res_48_45,wire_res_48_44,wire_res_48_43,wire_res_48_42,wire_res_48_41,
    wire_res_48_40,wire_res_48_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_24_lo = {wire_res_48_52,wire_res_48_51,wire_res_48_50,wire_res_48_49,wire_res_48_48,
    wire_res_48_47,wire_res_48_46,result_reg_r_24_lo_hi_hi_lo,result_reg_r_24_lo_hi_lo,result_reg_r_24_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_24_hi_lo_lo_lo = {wire_res_48_58,wire_res_48_57,wire_res_48_56,wire_res_48_55,wire_res_48_54,
    wire_res_48_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_24_hi_lo_lo = {wire_res_48_65,wire_res_48_64,wire_res_48_63,wire_res_48_62,wire_res_48_61,
    wire_res_48_60,wire_res_48_59,result_reg_r_24_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_24_hi_lo_hi_lo = {wire_res_48_71,wire_res_48_70,wire_res_48_69,wire_res_48_68,wire_res_48_67,
    wire_res_48_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_24_hi_lo = {wire_res_48_78,wire_res_48_77,wire_res_48_76,wire_res_48_75,wire_res_48_74,
    wire_res_48_73,wire_res_48_72,result_reg_r_24_hi_lo_hi_lo,result_reg_r_24_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_24_hi_hi_lo_lo = {wire_res_48_84,wire_res_48_83,wire_res_48_82,wire_res_48_81,wire_res_48_80,
    wire_res_48_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_24_hi_hi_lo = {wire_res_48_91,wire_res_48_90,wire_res_48_89,wire_res_48_88,wire_res_48_87,
    wire_res_48_86,wire_res_48_85,result_reg_r_24_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_24_hi_hi_hi_lo = {wire_res_48_98,wire_res_48_97,wire_res_48_96,wire_res_48_95,wire_res_48_94,
    wire_res_48_93,wire_res_48_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_24_hi = {wire_res_48_105,wire_res_48_104,wire_res_48_103,wire_res_48_102,wire_res_48_101,
    wire_res_48_100,wire_res_48_99,result_reg_r_24_hi_hi_hi_lo,result_reg_r_24_hi_hi_lo,result_reg_r_24_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_24_T = {result_reg_r_24_hi,result_reg_r_24_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [160:0] _a_aux_reg_w_25_T_2 = _GEN_1296 - _T_11336; // @[BinaryDesigns2.scala 225:48]
  wire [160:0] _GEN_100 = wire_res_49_55 ? _a_aux_reg_w_25_T_2 : {{55'd0}, a_aux_reg_r_24}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [159:0] _T_11338 = {b_aux_reg_r_24, 54'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_25 = _GEN_100[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [159:0] _GEN_1399 = {{54'd0}, a_aux_reg_w_25}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_50_54 = _GEN_1399 >= _T_11338; // @[BinaryDesigns2.scala 224:35]
  wire [159:0] _a_aux_reg_r_25_T_2 = _GEN_1399 - _T_11338; // @[BinaryDesigns2.scala 225:48]
  wire [159:0] _GEN_102 = wire_res_50_54 ? _a_aux_reg_r_25_T_2 : {{54'd0}, a_aux_reg_w_25}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_25_lo_lo_lo_lo = {wire_res_50_5,wire_res_50_4,wire_res_50_3,wire_res_50_2,wire_res_50_1,
    wire_res_50_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_25_lo_lo_lo = {wire_res_50_12,wire_res_50_11,wire_res_50_10,wire_res_50_9,wire_res_50_8,
    wire_res_50_7,wire_res_50_6,result_reg_r_25_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_25_lo_lo_hi_lo = {wire_res_50_18,wire_res_50_17,wire_res_50_16,wire_res_50_15,wire_res_50_14,
    wire_res_50_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_25_lo_lo = {wire_res_50_25,wire_res_50_24,wire_res_50_23,wire_res_50_22,wire_res_50_21,
    wire_res_50_20,wire_res_50_19,result_reg_r_25_lo_lo_hi_lo,result_reg_r_25_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_25_lo_hi_lo_lo = {wire_res_50_31,wire_res_50_30,wire_res_50_29,wire_res_50_28,wire_res_50_27,
    wire_res_50_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_25_lo_hi_lo = {wire_res_50_38,wire_res_50_37,wire_res_50_36,wire_res_50_35,wire_res_50_34,
    wire_res_50_33,wire_res_50_32,result_reg_r_25_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_25_lo_hi_hi_lo = {wire_res_50_45,wire_res_50_44,wire_res_50_43,wire_res_50_42,wire_res_50_41,
    wire_res_50_40,wire_res_50_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_25_lo = {wire_res_50_52,wire_res_50_51,wire_res_50_50,wire_res_50_49,wire_res_50_48,
    wire_res_50_47,wire_res_50_46,result_reg_r_25_lo_hi_hi_lo,result_reg_r_25_lo_hi_lo,result_reg_r_25_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_25_hi_lo_lo_lo = {wire_res_50_58,wire_res_50_57,wire_res_50_56,wire_res_50_55,wire_res_50_54,
    wire_res_50_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_25_hi_lo_lo = {wire_res_50_65,wire_res_50_64,wire_res_50_63,wire_res_50_62,wire_res_50_61,
    wire_res_50_60,wire_res_50_59,result_reg_r_25_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_25_hi_lo_hi_lo = {wire_res_50_71,wire_res_50_70,wire_res_50_69,wire_res_50_68,wire_res_50_67,
    wire_res_50_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_25_hi_lo = {wire_res_50_78,wire_res_50_77,wire_res_50_76,wire_res_50_75,wire_res_50_74,
    wire_res_50_73,wire_res_50_72,result_reg_r_25_hi_lo_hi_lo,result_reg_r_25_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_25_hi_hi_lo_lo = {wire_res_50_84,wire_res_50_83,wire_res_50_82,wire_res_50_81,wire_res_50_80,
    wire_res_50_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_25_hi_hi_lo = {wire_res_50_91,wire_res_50_90,wire_res_50_89,wire_res_50_88,wire_res_50_87,
    wire_res_50_86,wire_res_50_85,result_reg_r_25_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_25_hi_hi_hi_lo = {wire_res_50_98,wire_res_50_97,wire_res_50_96,wire_res_50_95,wire_res_50_94,
    wire_res_50_93,wire_res_50_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_25_hi = {wire_res_50_105,wire_res_50_104,wire_res_50_103,wire_res_50_102,wire_res_50_101,
    wire_res_50_100,wire_res_50_99,result_reg_r_25_hi_hi_hi_lo,result_reg_r_25_hi_hi_lo,result_reg_r_25_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_25_T = {result_reg_r_25_hi,result_reg_r_25_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [158:0] _a_aux_reg_w_26_T_2 = _GEN_1297 - _T_11340; // @[BinaryDesigns2.scala 225:48]
  wire [158:0] _GEN_104 = wire_res_51_53 ? _a_aux_reg_w_26_T_2 : {{53'd0}, a_aux_reg_r_25}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [157:0] _T_11342 = {b_aux_reg_r_25, 52'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_26 = _GEN_104[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [157:0] _GEN_1402 = {{52'd0}, a_aux_reg_w_26}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_52_52 = _GEN_1402 >= _T_11342; // @[BinaryDesigns2.scala 224:35]
  wire [157:0] _a_aux_reg_r_26_T_2 = _GEN_1402 - _T_11342; // @[BinaryDesigns2.scala 225:48]
  wire [157:0] _GEN_106 = wire_res_52_52 ? _a_aux_reg_r_26_T_2 : {{52'd0}, a_aux_reg_w_26}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_26_lo_lo_lo_lo = {wire_res_52_5,wire_res_52_4,wire_res_52_3,wire_res_52_2,wire_res_52_1,
    wire_res_52_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_26_lo_lo_lo = {wire_res_52_12,wire_res_52_11,wire_res_52_10,wire_res_52_9,wire_res_52_8,
    wire_res_52_7,wire_res_52_6,result_reg_r_26_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_26_lo_lo_hi_lo = {wire_res_52_18,wire_res_52_17,wire_res_52_16,wire_res_52_15,wire_res_52_14,
    wire_res_52_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_26_lo_lo = {wire_res_52_25,wire_res_52_24,wire_res_52_23,wire_res_52_22,wire_res_52_21,
    wire_res_52_20,wire_res_52_19,result_reg_r_26_lo_lo_hi_lo,result_reg_r_26_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_26_lo_hi_lo_lo = {wire_res_52_31,wire_res_52_30,wire_res_52_29,wire_res_52_28,wire_res_52_27,
    wire_res_52_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_26_lo_hi_lo = {wire_res_52_38,wire_res_52_37,wire_res_52_36,wire_res_52_35,wire_res_52_34,
    wire_res_52_33,wire_res_52_32,result_reg_r_26_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_26_lo_hi_hi_lo = {wire_res_52_45,wire_res_52_44,wire_res_52_43,wire_res_52_42,wire_res_52_41,
    wire_res_52_40,wire_res_52_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_26_lo = {wire_res_52_52,wire_res_52_51,wire_res_52_50,wire_res_52_49,wire_res_52_48,
    wire_res_52_47,wire_res_52_46,result_reg_r_26_lo_hi_hi_lo,result_reg_r_26_lo_hi_lo,result_reg_r_26_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_26_hi_lo_lo_lo = {wire_res_52_58,wire_res_52_57,wire_res_52_56,wire_res_52_55,wire_res_52_54,
    wire_res_52_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_26_hi_lo_lo = {wire_res_52_65,wire_res_52_64,wire_res_52_63,wire_res_52_62,wire_res_52_61,
    wire_res_52_60,wire_res_52_59,result_reg_r_26_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_26_hi_lo_hi_lo = {wire_res_52_71,wire_res_52_70,wire_res_52_69,wire_res_52_68,wire_res_52_67,
    wire_res_52_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_26_hi_lo = {wire_res_52_78,wire_res_52_77,wire_res_52_76,wire_res_52_75,wire_res_52_74,
    wire_res_52_73,wire_res_52_72,result_reg_r_26_hi_lo_hi_lo,result_reg_r_26_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_26_hi_hi_lo_lo = {wire_res_52_84,wire_res_52_83,wire_res_52_82,wire_res_52_81,wire_res_52_80,
    wire_res_52_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_26_hi_hi_lo = {wire_res_52_91,wire_res_52_90,wire_res_52_89,wire_res_52_88,wire_res_52_87,
    wire_res_52_86,wire_res_52_85,result_reg_r_26_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_26_hi_hi_hi_lo = {wire_res_52_98,wire_res_52_97,wire_res_52_96,wire_res_52_95,wire_res_52_94,
    wire_res_52_93,wire_res_52_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_26_hi = {wire_res_52_105,wire_res_52_104,wire_res_52_103,wire_res_52_102,wire_res_52_101,
    wire_res_52_100,wire_res_52_99,result_reg_r_26_hi_hi_hi_lo,result_reg_r_26_hi_hi_lo,result_reg_r_26_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_26_T = {result_reg_r_26_hi,result_reg_r_26_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [156:0] _a_aux_reg_w_27_T_2 = _GEN_1298 - _T_11344; // @[BinaryDesigns2.scala 225:48]
  wire [156:0] _GEN_108 = wire_res_53_51 ? _a_aux_reg_w_27_T_2 : {{51'd0}, a_aux_reg_r_26}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [155:0] _T_11346 = {b_aux_reg_r_26, 50'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_27 = _GEN_108[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [155:0] _GEN_1405 = {{50'd0}, a_aux_reg_w_27}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_54_50 = _GEN_1405 >= _T_11346; // @[BinaryDesigns2.scala 224:35]
  wire [155:0] _a_aux_reg_r_27_T_2 = _GEN_1405 - _T_11346; // @[BinaryDesigns2.scala 225:48]
  wire [155:0] _GEN_110 = wire_res_54_50 ? _a_aux_reg_r_27_T_2 : {{50'd0}, a_aux_reg_w_27}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_27_lo_lo_lo_lo = {wire_res_54_5,wire_res_54_4,wire_res_54_3,wire_res_54_2,wire_res_54_1,
    wire_res_54_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_27_lo_lo_lo = {wire_res_54_12,wire_res_54_11,wire_res_54_10,wire_res_54_9,wire_res_54_8,
    wire_res_54_7,wire_res_54_6,result_reg_r_27_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_27_lo_lo_hi_lo = {wire_res_54_18,wire_res_54_17,wire_res_54_16,wire_res_54_15,wire_res_54_14,
    wire_res_54_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_27_lo_lo = {wire_res_54_25,wire_res_54_24,wire_res_54_23,wire_res_54_22,wire_res_54_21,
    wire_res_54_20,wire_res_54_19,result_reg_r_27_lo_lo_hi_lo,result_reg_r_27_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_27_lo_hi_lo_lo = {wire_res_54_31,wire_res_54_30,wire_res_54_29,wire_res_54_28,wire_res_54_27,
    wire_res_54_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_27_lo_hi_lo = {wire_res_54_38,wire_res_54_37,wire_res_54_36,wire_res_54_35,wire_res_54_34,
    wire_res_54_33,wire_res_54_32,result_reg_r_27_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_27_lo_hi_hi_lo = {wire_res_54_45,wire_res_54_44,wire_res_54_43,wire_res_54_42,wire_res_54_41,
    wire_res_54_40,wire_res_54_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_27_lo = {wire_res_54_52,wire_res_54_51,wire_res_54_50,wire_res_54_49,wire_res_54_48,
    wire_res_54_47,wire_res_54_46,result_reg_r_27_lo_hi_hi_lo,result_reg_r_27_lo_hi_lo,result_reg_r_27_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_27_hi_lo_lo_lo = {wire_res_54_58,wire_res_54_57,wire_res_54_56,wire_res_54_55,wire_res_54_54,
    wire_res_54_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_27_hi_lo_lo = {wire_res_54_65,wire_res_54_64,wire_res_54_63,wire_res_54_62,wire_res_54_61,
    wire_res_54_60,wire_res_54_59,result_reg_r_27_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_27_hi_lo_hi_lo = {wire_res_54_71,wire_res_54_70,wire_res_54_69,wire_res_54_68,wire_res_54_67,
    wire_res_54_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_27_hi_lo = {wire_res_54_78,wire_res_54_77,wire_res_54_76,wire_res_54_75,wire_res_54_74,
    wire_res_54_73,wire_res_54_72,result_reg_r_27_hi_lo_hi_lo,result_reg_r_27_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_27_hi_hi_lo_lo = {wire_res_54_84,wire_res_54_83,wire_res_54_82,wire_res_54_81,wire_res_54_80,
    wire_res_54_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_27_hi_hi_lo = {wire_res_54_91,wire_res_54_90,wire_res_54_89,wire_res_54_88,wire_res_54_87,
    wire_res_54_86,wire_res_54_85,result_reg_r_27_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_27_hi_hi_hi_lo = {wire_res_54_98,wire_res_54_97,wire_res_54_96,wire_res_54_95,wire_res_54_94,
    wire_res_54_93,wire_res_54_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_27_hi = {wire_res_54_105,wire_res_54_104,wire_res_54_103,wire_res_54_102,wire_res_54_101,
    wire_res_54_100,wire_res_54_99,result_reg_r_27_hi_hi_hi_lo,result_reg_r_27_hi_hi_lo,result_reg_r_27_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_27_T = {result_reg_r_27_hi,result_reg_r_27_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [154:0] _a_aux_reg_w_28_T_2 = _GEN_1299 - _T_11348; // @[BinaryDesigns2.scala 225:48]
  wire [154:0] _GEN_112 = wire_res_55_49 ? _a_aux_reg_w_28_T_2 : {{49'd0}, a_aux_reg_r_27}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [153:0] _T_11350 = {b_aux_reg_r_27, 48'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_28 = _GEN_112[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [153:0] _GEN_1408 = {{48'd0}, a_aux_reg_w_28}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_56_48 = _GEN_1408 >= _T_11350; // @[BinaryDesigns2.scala 224:35]
  wire [153:0] _a_aux_reg_r_28_T_2 = _GEN_1408 - _T_11350; // @[BinaryDesigns2.scala 225:48]
  wire [153:0] _GEN_114 = wire_res_56_48 ? _a_aux_reg_r_28_T_2 : {{48'd0}, a_aux_reg_w_28}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_28_lo_lo_lo_lo = {wire_res_56_5,wire_res_56_4,wire_res_56_3,wire_res_56_2,wire_res_56_1,
    wire_res_56_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_28_lo_lo_lo = {wire_res_56_12,wire_res_56_11,wire_res_56_10,wire_res_56_9,wire_res_56_8,
    wire_res_56_7,wire_res_56_6,result_reg_r_28_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_28_lo_lo_hi_lo = {wire_res_56_18,wire_res_56_17,wire_res_56_16,wire_res_56_15,wire_res_56_14,
    wire_res_56_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_28_lo_lo = {wire_res_56_25,wire_res_56_24,wire_res_56_23,wire_res_56_22,wire_res_56_21,
    wire_res_56_20,wire_res_56_19,result_reg_r_28_lo_lo_hi_lo,result_reg_r_28_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_28_lo_hi_lo_lo = {wire_res_56_31,wire_res_56_30,wire_res_56_29,wire_res_56_28,wire_res_56_27,
    wire_res_56_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_28_lo_hi_lo = {wire_res_56_38,wire_res_56_37,wire_res_56_36,wire_res_56_35,wire_res_56_34,
    wire_res_56_33,wire_res_56_32,result_reg_r_28_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_28_lo_hi_hi_lo = {wire_res_56_45,wire_res_56_44,wire_res_56_43,wire_res_56_42,wire_res_56_41,
    wire_res_56_40,wire_res_56_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_28_lo = {wire_res_56_52,wire_res_56_51,wire_res_56_50,wire_res_56_49,wire_res_56_48,
    wire_res_56_47,wire_res_56_46,result_reg_r_28_lo_hi_hi_lo,result_reg_r_28_lo_hi_lo,result_reg_r_28_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_28_hi_lo_lo_lo = {wire_res_56_58,wire_res_56_57,wire_res_56_56,wire_res_56_55,wire_res_56_54,
    wire_res_56_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_28_hi_lo_lo = {wire_res_56_65,wire_res_56_64,wire_res_56_63,wire_res_56_62,wire_res_56_61,
    wire_res_56_60,wire_res_56_59,result_reg_r_28_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_28_hi_lo_hi_lo = {wire_res_56_71,wire_res_56_70,wire_res_56_69,wire_res_56_68,wire_res_56_67,
    wire_res_56_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_28_hi_lo = {wire_res_56_78,wire_res_56_77,wire_res_56_76,wire_res_56_75,wire_res_56_74,
    wire_res_56_73,wire_res_56_72,result_reg_r_28_hi_lo_hi_lo,result_reg_r_28_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_28_hi_hi_lo_lo = {wire_res_56_84,wire_res_56_83,wire_res_56_82,wire_res_56_81,wire_res_56_80,
    wire_res_56_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_28_hi_hi_lo = {wire_res_56_91,wire_res_56_90,wire_res_56_89,wire_res_56_88,wire_res_56_87,
    wire_res_56_86,wire_res_56_85,result_reg_r_28_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_28_hi_hi_hi_lo = {wire_res_56_98,wire_res_56_97,wire_res_56_96,wire_res_56_95,wire_res_56_94,
    wire_res_56_93,wire_res_56_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_28_hi = {wire_res_56_105,wire_res_56_104,wire_res_56_103,wire_res_56_102,wire_res_56_101,
    wire_res_56_100,wire_res_56_99,result_reg_r_28_hi_hi_hi_lo,result_reg_r_28_hi_hi_lo,result_reg_r_28_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_28_T = {result_reg_r_28_hi,result_reg_r_28_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [152:0] _a_aux_reg_w_29_T_2 = _GEN_1300 - _T_11352; // @[BinaryDesigns2.scala 225:48]
  wire [152:0] _GEN_116 = wire_res_57_47 ? _a_aux_reg_w_29_T_2 : {{47'd0}, a_aux_reg_r_28}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [151:0] _T_11354 = {b_aux_reg_r_28, 46'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_29 = _GEN_116[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [151:0] _GEN_1411 = {{46'd0}, a_aux_reg_w_29}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_58_46 = _GEN_1411 >= _T_11354; // @[BinaryDesigns2.scala 224:35]
  wire [151:0] _a_aux_reg_r_29_T_2 = _GEN_1411 - _T_11354; // @[BinaryDesigns2.scala 225:48]
  wire [151:0] _GEN_118 = wire_res_58_46 ? _a_aux_reg_r_29_T_2 : {{46'd0}, a_aux_reg_w_29}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_29_lo_lo_lo_lo = {wire_res_58_5,wire_res_58_4,wire_res_58_3,wire_res_58_2,wire_res_58_1,
    wire_res_58_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_29_lo_lo_lo = {wire_res_58_12,wire_res_58_11,wire_res_58_10,wire_res_58_9,wire_res_58_8,
    wire_res_58_7,wire_res_58_6,result_reg_r_29_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_29_lo_lo_hi_lo = {wire_res_58_18,wire_res_58_17,wire_res_58_16,wire_res_58_15,wire_res_58_14,
    wire_res_58_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_29_lo_lo = {wire_res_58_25,wire_res_58_24,wire_res_58_23,wire_res_58_22,wire_res_58_21,
    wire_res_58_20,wire_res_58_19,result_reg_r_29_lo_lo_hi_lo,result_reg_r_29_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_29_lo_hi_lo_lo = {wire_res_58_31,wire_res_58_30,wire_res_58_29,wire_res_58_28,wire_res_58_27,
    wire_res_58_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_29_lo_hi_lo = {wire_res_58_38,wire_res_58_37,wire_res_58_36,wire_res_58_35,wire_res_58_34,
    wire_res_58_33,wire_res_58_32,result_reg_r_29_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_29_lo_hi_hi_lo = {wire_res_58_45,wire_res_58_44,wire_res_58_43,wire_res_58_42,wire_res_58_41,
    wire_res_58_40,wire_res_58_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_29_lo = {wire_res_58_52,wire_res_58_51,wire_res_58_50,wire_res_58_49,wire_res_58_48,
    wire_res_58_47,wire_res_58_46,result_reg_r_29_lo_hi_hi_lo,result_reg_r_29_lo_hi_lo,result_reg_r_29_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_29_hi_lo_lo_lo = {wire_res_58_58,wire_res_58_57,wire_res_58_56,wire_res_58_55,wire_res_58_54,
    wire_res_58_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_29_hi_lo_lo = {wire_res_58_65,wire_res_58_64,wire_res_58_63,wire_res_58_62,wire_res_58_61,
    wire_res_58_60,wire_res_58_59,result_reg_r_29_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_29_hi_lo_hi_lo = {wire_res_58_71,wire_res_58_70,wire_res_58_69,wire_res_58_68,wire_res_58_67,
    wire_res_58_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_29_hi_lo = {wire_res_58_78,wire_res_58_77,wire_res_58_76,wire_res_58_75,wire_res_58_74,
    wire_res_58_73,wire_res_58_72,result_reg_r_29_hi_lo_hi_lo,result_reg_r_29_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_29_hi_hi_lo_lo = {wire_res_58_84,wire_res_58_83,wire_res_58_82,wire_res_58_81,wire_res_58_80,
    wire_res_58_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_29_hi_hi_lo = {wire_res_58_91,wire_res_58_90,wire_res_58_89,wire_res_58_88,wire_res_58_87,
    wire_res_58_86,wire_res_58_85,result_reg_r_29_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_29_hi_hi_hi_lo = {wire_res_58_98,wire_res_58_97,wire_res_58_96,wire_res_58_95,wire_res_58_94,
    wire_res_58_93,wire_res_58_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_29_hi = {wire_res_58_105,wire_res_58_104,wire_res_58_103,wire_res_58_102,wire_res_58_101,
    wire_res_58_100,wire_res_58_99,result_reg_r_29_hi_hi_hi_lo,result_reg_r_29_hi_hi_lo,result_reg_r_29_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_29_T = {result_reg_r_29_hi,result_reg_r_29_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [150:0] _a_aux_reg_w_30_T_2 = _GEN_1301 - _T_11356; // @[BinaryDesigns2.scala 225:48]
  wire [150:0] _GEN_120 = wire_res_59_45 ? _a_aux_reg_w_30_T_2 : {{45'd0}, a_aux_reg_r_29}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [149:0] _T_11358 = {b_aux_reg_r_29, 44'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_30 = _GEN_120[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [149:0] _GEN_1414 = {{44'd0}, a_aux_reg_w_30}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_60_44 = _GEN_1414 >= _T_11358; // @[BinaryDesigns2.scala 224:35]
  wire [149:0] _a_aux_reg_r_30_T_2 = _GEN_1414 - _T_11358; // @[BinaryDesigns2.scala 225:48]
  wire [149:0] _GEN_122 = wire_res_60_44 ? _a_aux_reg_r_30_T_2 : {{44'd0}, a_aux_reg_w_30}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_30_lo_lo_lo_lo = {wire_res_60_5,wire_res_60_4,wire_res_60_3,wire_res_60_2,wire_res_60_1,
    wire_res_60_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_30_lo_lo_lo = {wire_res_60_12,wire_res_60_11,wire_res_60_10,wire_res_60_9,wire_res_60_8,
    wire_res_60_7,wire_res_60_6,result_reg_r_30_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_30_lo_lo_hi_lo = {wire_res_60_18,wire_res_60_17,wire_res_60_16,wire_res_60_15,wire_res_60_14,
    wire_res_60_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_30_lo_lo = {wire_res_60_25,wire_res_60_24,wire_res_60_23,wire_res_60_22,wire_res_60_21,
    wire_res_60_20,wire_res_60_19,result_reg_r_30_lo_lo_hi_lo,result_reg_r_30_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_30_lo_hi_lo_lo = {wire_res_60_31,wire_res_60_30,wire_res_60_29,wire_res_60_28,wire_res_60_27,
    wire_res_60_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_30_lo_hi_lo = {wire_res_60_38,wire_res_60_37,wire_res_60_36,wire_res_60_35,wire_res_60_34,
    wire_res_60_33,wire_res_60_32,result_reg_r_30_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_30_lo_hi_hi_lo = {wire_res_60_45,wire_res_60_44,wire_res_60_43,wire_res_60_42,wire_res_60_41,
    wire_res_60_40,wire_res_60_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_30_lo = {wire_res_60_52,wire_res_60_51,wire_res_60_50,wire_res_60_49,wire_res_60_48,
    wire_res_60_47,wire_res_60_46,result_reg_r_30_lo_hi_hi_lo,result_reg_r_30_lo_hi_lo,result_reg_r_30_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_30_hi_lo_lo_lo = {wire_res_60_58,wire_res_60_57,wire_res_60_56,wire_res_60_55,wire_res_60_54,
    wire_res_60_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_30_hi_lo_lo = {wire_res_60_65,wire_res_60_64,wire_res_60_63,wire_res_60_62,wire_res_60_61,
    wire_res_60_60,wire_res_60_59,result_reg_r_30_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_30_hi_lo_hi_lo = {wire_res_60_71,wire_res_60_70,wire_res_60_69,wire_res_60_68,wire_res_60_67,
    wire_res_60_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_30_hi_lo = {wire_res_60_78,wire_res_60_77,wire_res_60_76,wire_res_60_75,wire_res_60_74,
    wire_res_60_73,wire_res_60_72,result_reg_r_30_hi_lo_hi_lo,result_reg_r_30_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_30_hi_hi_lo_lo = {wire_res_60_84,wire_res_60_83,wire_res_60_82,wire_res_60_81,wire_res_60_80,
    wire_res_60_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_30_hi_hi_lo = {wire_res_60_91,wire_res_60_90,wire_res_60_89,wire_res_60_88,wire_res_60_87,
    wire_res_60_86,wire_res_60_85,result_reg_r_30_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_30_hi_hi_hi_lo = {wire_res_60_98,wire_res_60_97,wire_res_60_96,wire_res_60_95,wire_res_60_94,
    wire_res_60_93,wire_res_60_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_30_hi = {wire_res_60_105,wire_res_60_104,wire_res_60_103,wire_res_60_102,wire_res_60_101,
    wire_res_60_100,wire_res_60_99,result_reg_r_30_hi_hi_hi_lo,result_reg_r_30_hi_hi_lo,result_reg_r_30_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_30_T = {result_reg_r_30_hi,result_reg_r_30_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [148:0] _a_aux_reg_w_31_T_2 = _GEN_1302 - _T_11360; // @[BinaryDesigns2.scala 225:48]
  wire [148:0] _GEN_124 = wire_res_61_43 ? _a_aux_reg_w_31_T_2 : {{43'd0}, a_aux_reg_r_30}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [147:0] _T_11362 = {b_aux_reg_r_30, 42'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_31 = _GEN_124[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [147:0] _GEN_1417 = {{42'd0}, a_aux_reg_w_31}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_62_42 = _GEN_1417 >= _T_11362; // @[BinaryDesigns2.scala 224:35]
  wire [147:0] _a_aux_reg_r_31_T_2 = _GEN_1417 - _T_11362; // @[BinaryDesigns2.scala 225:48]
  wire [147:0] _GEN_126 = wire_res_62_42 ? _a_aux_reg_r_31_T_2 : {{42'd0}, a_aux_reg_w_31}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_31_lo_lo_lo_lo = {wire_res_62_5,wire_res_62_4,wire_res_62_3,wire_res_62_2,wire_res_62_1,
    wire_res_62_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_31_lo_lo_lo = {wire_res_62_12,wire_res_62_11,wire_res_62_10,wire_res_62_9,wire_res_62_8,
    wire_res_62_7,wire_res_62_6,result_reg_r_31_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_31_lo_lo_hi_lo = {wire_res_62_18,wire_res_62_17,wire_res_62_16,wire_res_62_15,wire_res_62_14,
    wire_res_62_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_31_lo_lo = {wire_res_62_25,wire_res_62_24,wire_res_62_23,wire_res_62_22,wire_res_62_21,
    wire_res_62_20,wire_res_62_19,result_reg_r_31_lo_lo_hi_lo,result_reg_r_31_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_31_lo_hi_lo_lo = {wire_res_62_31,wire_res_62_30,wire_res_62_29,wire_res_62_28,wire_res_62_27,
    wire_res_62_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_31_lo_hi_lo = {wire_res_62_38,wire_res_62_37,wire_res_62_36,wire_res_62_35,wire_res_62_34,
    wire_res_62_33,wire_res_62_32,result_reg_r_31_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_31_lo_hi_hi_lo = {wire_res_62_45,wire_res_62_44,wire_res_62_43,wire_res_62_42,wire_res_62_41,
    wire_res_62_40,wire_res_62_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_31_lo = {wire_res_62_52,wire_res_62_51,wire_res_62_50,wire_res_62_49,wire_res_62_48,
    wire_res_62_47,wire_res_62_46,result_reg_r_31_lo_hi_hi_lo,result_reg_r_31_lo_hi_lo,result_reg_r_31_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_31_hi_lo_lo_lo = {wire_res_62_58,wire_res_62_57,wire_res_62_56,wire_res_62_55,wire_res_62_54,
    wire_res_62_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_31_hi_lo_lo = {wire_res_62_65,wire_res_62_64,wire_res_62_63,wire_res_62_62,wire_res_62_61,
    wire_res_62_60,wire_res_62_59,result_reg_r_31_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_31_hi_lo_hi_lo = {wire_res_62_71,wire_res_62_70,wire_res_62_69,wire_res_62_68,wire_res_62_67,
    wire_res_62_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_31_hi_lo = {wire_res_62_78,wire_res_62_77,wire_res_62_76,wire_res_62_75,wire_res_62_74,
    wire_res_62_73,wire_res_62_72,result_reg_r_31_hi_lo_hi_lo,result_reg_r_31_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_31_hi_hi_lo_lo = {wire_res_62_84,wire_res_62_83,wire_res_62_82,wire_res_62_81,wire_res_62_80,
    wire_res_62_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_31_hi_hi_lo = {wire_res_62_91,wire_res_62_90,wire_res_62_89,wire_res_62_88,wire_res_62_87,
    wire_res_62_86,wire_res_62_85,result_reg_r_31_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_31_hi_hi_hi_lo = {wire_res_62_98,wire_res_62_97,wire_res_62_96,wire_res_62_95,wire_res_62_94,
    wire_res_62_93,wire_res_62_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_31_hi = {wire_res_62_105,wire_res_62_104,wire_res_62_103,wire_res_62_102,wire_res_62_101,
    wire_res_62_100,wire_res_62_99,result_reg_r_31_hi_hi_hi_lo,result_reg_r_31_hi_hi_lo,result_reg_r_31_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_31_T = {result_reg_r_31_hi,result_reg_r_31_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [146:0] _a_aux_reg_w_32_T_2 = _GEN_1303 - _T_11364; // @[BinaryDesigns2.scala 225:48]
  wire [146:0] _GEN_128 = wire_res_63_41 ? _a_aux_reg_w_32_T_2 : {{41'd0}, a_aux_reg_r_31}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [145:0] _T_11366 = {b_aux_reg_r_31, 40'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_32 = _GEN_128[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [145:0] _GEN_1420 = {{40'd0}, a_aux_reg_w_32}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_64_40 = _GEN_1420 >= _T_11366; // @[BinaryDesigns2.scala 224:35]
  wire [145:0] _a_aux_reg_r_32_T_2 = _GEN_1420 - _T_11366; // @[BinaryDesigns2.scala 225:48]
  wire [145:0] _GEN_130 = wire_res_64_40 ? _a_aux_reg_r_32_T_2 : {{40'd0}, a_aux_reg_w_32}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_32_lo_lo_lo_lo = {wire_res_64_5,wire_res_64_4,wire_res_64_3,wire_res_64_2,wire_res_64_1,
    wire_res_64_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_32_lo_lo_lo = {wire_res_64_12,wire_res_64_11,wire_res_64_10,wire_res_64_9,wire_res_64_8,
    wire_res_64_7,wire_res_64_6,result_reg_r_32_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_32_lo_lo_hi_lo = {wire_res_64_18,wire_res_64_17,wire_res_64_16,wire_res_64_15,wire_res_64_14,
    wire_res_64_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_32_lo_lo = {wire_res_64_25,wire_res_64_24,wire_res_64_23,wire_res_64_22,wire_res_64_21,
    wire_res_64_20,wire_res_64_19,result_reg_r_32_lo_lo_hi_lo,result_reg_r_32_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_32_lo_hi_lo_lo = {wire_res_64_31,wire_res_64_30,wire_res_64_29,wire_res_64_28,wire_res_64_27,
    wire_res_64_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_32_lo_hi_lo = {wire_res_64_38,wire_res_64_37,wire_res_64_36,wire_res_64_35,wire_res_64_34,
    wire_res_64_33,wire_res_64_32,result_reg_r_32_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_32_lo_hi_hi_lo = {wire_res_64_45,wire_res_64_44,wire_res_64_43,wire_res_64_42,wire_res_64_41,
    wire_res_64_40,wire_res_64_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_32_lo = {wire_res_64_52,wire_res_64_51,wire_res_64_50,wire_res_64_49,wire_res_64_48,
    wire_res_64_47,wire_res_64_46,result_reg_r_32_lo_hi_hi_lo,result_reg_r_32_lo_hi_lo,result_reg_r_32_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_32_hi_lo_lo_lo = {wire_res_64_58,wire_res_64_57,wire_res_64_56,wire_res_64_55,wire_res_64_54,
    wire_res_64_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_32_hi_lo_lo = {wire_res_64_65,wire_res_64_64,wire_res_64_63,wire_res_64_62,wire_res_64_61,
    wire_res_64_60,wire_res_64_59,result_reg_r_32_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_32_hi_lo_hi_lo = {wire_res_64_71,wire_res_64_70,wire_res_64_69,wire_res_64_68,wire_res_64_67,
    wire_res_64_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_32_hi_lo = {wire_res_64_78,wire_res_64_77,wire_res_64_76,wire_res_64_75,wire_res_64_74,
    wire_res_64_73,wire_res_64_72,result_reg_r_32_hi_lo_hi_lo,result_reg_r_32_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_32_hi_hi_lo_lo = {wire_res_64_84,wire_res_64_83,wire_res_64_82,wire_res_64_81,wire_res_64_80,
    wire_res_64_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_32_hi_hi_lo = {wire_res_64_91,wire_res_64_90,wire_res_64_89,wire_res_64_88,wire_res_64_87,
    wire_res_64_86,wire_res_64_85,result_reg_r_32_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_32_hi_hi_hi_lo = {wire_res_64_98,wire_res_64_97,wire_res_64_96,wire_res_64_95,wire_res_64_94,
    wire_res_64_93,wire_res_64_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_32_hi = {wire_res_64_105,wire_res_64_104,wire_res_64_103,wire_res_64_102,wire_res_64_101,
    wire_res_64_100,wire_res_64_99,result_reg_r_32_hi_hi_hi_lo,result_reg_r_32_hi_hi_lo,result_reg_r_32_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_32_T = {result_reg_r_32_hi,result_reg_r_32_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [144:0] _a_aux_reg_w_33_T_2 = _GEN_1304 - _T_11368; // @[BinaryDesigns2.scala 225:48]
  wire [144:0] _GEN_132 = wire_res_65_39 ? _a_aux_reg_w_33_T_2 : {{39'd0}, a_aux_reg_r_32}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [143:0] _T_11370 = {b_aux_reg_r_32, 38'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_33 = _GEN_132[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [143:0] _GEN_1423 = {{38'd0}, a_aux_reg_w_33}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_66_38 = _GEN_1423 >= _T_11370; // @[BinaryDesigns2.scala 224:35]
  wire [143:0] _a_aux_reg_r_33_T_2 = _GEN_1423 - _T_11370; // @[BinaryDesigns2.scala 225:48]
  wire [143:0] _GEN_134 = wire_res_66_38 ? _a_aux_reg_r_33_T_2 : {{38'd0}, a_aux_reg_w_33}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_33_lo_lo_lo_lo = {wire_res_66_5,wire_res_66_4,wire_res_66_3,wire_res_66_2,wire_res_66_1,
    wire_res_66_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_33_lo_lo_lo = {wire_res_66_12,wire_res_66_11,wire_res_66_10,wire_res_66_9,wire_res_66_8,
    wire_res_66_7,wire_res_66_6,result_reg_r_33_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_33_lo_lo_hi_lo = {wire_res_66_18,wire_res_66_17,wire_res_66_16,wire_res_66_15,wire_res_66_14,
    wire_res_66_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_33_lo_lo = {wire_res_66_25,wire_res_66_24,wire_res_66_23,wire_res_66_22,wire_res_66_21,
    wire_res_66_20,wire_res_66_19,result_reg_r_33_lo_lo_hi_lo,result_reg_r_33_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_33_lo_hi_lo_lo = {wire_res_66_31,wire_res_66_30,wire_res_66_29,wire_res_66_28,wire_res_66_27,
    wire_res_66_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_33_lo_hi_lo = {wire_res_66_38,wire_res_66_37,wire_res_66_36,wire_res_66_35,wire_res_66_34,
    wire_res_66_33,wire_res_66_32,result_reg_r_33_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_33_lo_hi_hi_lo = {wire_res_66_45,wire_res_66_44,wire_res_66_43,wire_res_66_42,wire_res_66_41,
    wire_res_66_40,wire_res_66_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_33_lo = {wire_res_66_52,wire_res_66_51,wire_res_66_50,wire_res_66_49,wire_res_66_48,
    wire_res_66_47,wire_res_66_46,result_reg_r_33_lo_hi_hi_lo,result_reg_r_33_lo_hi_lo,result_reg_r_33_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_33_hi_lo_lo_lo = {wire_res_66_58,wire_res_66_57,wire_res_66_56,wire_res_66_55,wire_res_66_54,
    wire_res_66_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_33_hi_lo_lo = {wire_res_66_65,wire_res_66_64,wire_res_66_63,wire_res_66_62,wire_res_66_61,
    wire_res_66_60,wire_res_66_59,result_reg_r_33_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_33_hi_lo_hi_lo = {wire_res_66_71,wire_res_66_70,wire_res_66_69,wire_res_66_68,wire_res_66_67,
    wire_res_66_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_33_hi_lo = {wire_res_66_78,wire_res_66_77,wire_res_66_76,wire_res_66_75,wire_res_66_74,
    wire_res_66_73,wire_res_66_72,result_reg_r_33_hi_lo_hi_lo,result_reg_r_33_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_33_hi_hi_lo_lo = {wire_res_66_84,wire_res_66_83,wire_res_66_82,wire_res_66_81,wire_res_66_80,
    wire_res_66_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_33_hi_hi_lo = {wire_res_66_91,wire_res_66_90,wire_res_66_89,wire_res_66_88,wire_res_66_87,
    wire_res_66_86,wire_res_66_85,result_reg_r_33_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_33_hi_hi_hi_lo = {wire_res_66_98,wire_res_66_97,wire_res_66_96,wire_res_66_95,wire_res_66_94,
    wire_res_66_93,wire_res_66_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_33_hi = {wire_res_66_105,wire_res_66_104,wire_res_66_103,wire_res_66_102,wire_res_66_101,
    wire_res_66_100,wire_res_66_99,result_reg_r_33_hi_hi_hi_lo,result_reg_r_33_hi_hi_lo,result_reg_r_33_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_33_T = {result_reg_r_33_hi,result_reg_r_33_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [142:0] _a_aux_reg_w_34_T_2 = _GEN_1305 - _T_11372; // @[BinaryDesigns2.scala 225:48]
  wire [142:0] _GEN_136 = wire_res_67_37 ? _a_aux_reg_w_34_T_2 : {{37'd0}, a_aux_reg_r_33}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [141:0] _T_11374 = {b_aux_reg_r_33, 36'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_34 = _GEN_136[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [141:0] _GEN_1426 = {{36'd0}, a_aux_reg_w_34}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_68_36 = _GEN_1426 >= _T_11374; // @[BinaryDesigns2.scala 224:35]
  wire [141:0] _a_aux_reg_r_34_T_2 = _GEN_1426 - _T_11374; // @[BinaryDesigns2.scala 225:48]
  wire [141:0] _GEN_138 = wire_res_68_36 ? _a_aux_reg_r_34_T_2 : {{36'd0}, a_aux_reg_w_34}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_34_lo_lo_lo_lo = {wire_res_68_5,wire_res_68_4,wire_res_68_3,wire_res_68_2,wire_res_68_1,
    wire_res_68_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_34_lo_lo_lo = {wire_res_68_12,wire_res_68_11,wire_res_68_10,wire_res_68_9,wire_res_68_8,
    wire_res_68_7,wire_res_68_6,result_reg_r_34_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_34_lo_lo_hi_lo = {wire_res_68_18,wire_res_68_17,wire_res_68_16,wire_res_68_15,wire_res_68_14,
    wire_res_68_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_34_lo_lo = {wire_res_68_25,wire_res_68_24,wire_res_68_23,wire_res_68_22,wire_res_68_21,
    wire_res_68_20,wire_res_68_19,result_reg_r_34_lo_lo_hi_lo,result_reg_r_34_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_34_lo_hi_lo_lo = {wire_res_68_31,wire_res_68_30,wire_res_68_29,wire_res_68_28,wire_res_68_27,
    wire_res_68_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_34_lo_hi_lo = {wire_res_68_38,wire_res_68_37,wire_res_68_36,wire_res_68_35,wire_res_68_34,
    wire_res_68_33,wire_res_68_32,result_reg_r_34_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_34_lo_hi_hi_lo = {wire_res_68_45,wire_res_68_44,wire_res_68_43,wire_res_68_42,wire_res_68_41,
    wire_res_68_40,wire_res_68_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_34_lo = {wire_res_68_52,wire_res_68_51,wire_res_68_50,wire_res_68_49,wire_res_68_48,
    wire_res_68_47,wire_res_68_46,result_reg_r_34_lo_hi_hi_lo,result_reg_r_34_lo_hi_lo,result_reg_r_34_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_34_hi_lo_lo_lo = {wire_res_68_58,wire_res_68_57,wire_res_68_56,wire_res_68_55,wire_res_68_54,
    wire_res_68_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_34_hi_lo_lo = {wire_res_68_65,wire_res_68_64,wire_res_68_63,wire_res_68_62,wire_res_68_61,
    wire_res_68_60,wire_res_68_59,result_reg_r_34_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_34_hi_lo_hi_lo = {wire_res_68_71,wire_res_68_70,wire_res_68_69,wire_res_68_68,wire_res_68_67,
    wire_res_68_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_34_hi_lo = {wire_res_68_78,wire_res_68_77,wire_res_68_76,wire_res_68_75,wire_res_68_74,
    wire_res_68_73,wire_res_68_72,result_reg_r_34_hi_lo_hi_lo,result_reg_r_34_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_34_hi_hi_lo_lo = {wire_res_68_84,wire_res_68_83,wire_res_68_82,wire_res_68_81,wire_res_68_80,
    wire_res_68_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_34_hi_hi_lo = {wire_res_68_91,wire_res_68_90,wire_res_68_89,wire_res_68_88,wire_res_68_87,
    wire_res_68_86,wire_res_68_85,result_reg_r_34_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_34_hi_hi_hi_lo = {wire_res_68_98,wire_res_68_97,wire_res_68_96,wire_res_68_95,wire_res_68_94,
    wire_res_68_93,wire_res_68_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_34_hi = {wire_res_68_105,wire_res_68_104,wire_res_68_103,wire_res_68_102,wire_res_68_101,
    wire_res_68_100,wire_res_68_99,result_reg_r_34_hi_hi_hi_lo,result_reg_r_34_hi_hi_lo,result_reg_r_34_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_34_T = {result_reg_r_34_hi,result_reg_r_34_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [140:0] _a_aux_reg_w_35_T_2 = _GEN_1306 - _T_11376; // @[BinaryDesigns2.scala 225:48]
  wire [140:0] _GEN_140 = wire_res_69_35 ? _a_aux_reg_w_35_T_2 : {{35'd0}, a_aux_reg_r_34}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [139:0] _T_11378 = {b_aux_reg_r_34, 34'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_35 = _GEN_140[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [139:0] _GEN_1429 = {{34'd0}, a_aux_reg_w_35}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_70_34 = _GEN_1429 >= _T_11378; // @[BinaryDesigns2.scala 224:35]
  wire [139:0] _a_aux_reg_r_35_T_2 = _GEN_1429 - _T_11378; // @[BinaryDesigns2.scala 225:48]
  wire [139:0] _GEN_142 = wire_res_70_34 ? _a_aux_reg_r_35_T_2 : {{34'd0}, a_aux_reg_w_35}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_35_lo_lo_lo_lo = {wire_res_70_5,wire_res_70_4,wire_res_70_3,wire_res_70_2,wire_res_70_1,
    wire_res_70_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_35_lo_lo_lo = {wire_res_70_12,wire_res_70_11,wire_res_70_10,wire_res_70_9,wire_res_70_8,
    wire_res_70_7,wire_res_70_6,result_reg_r_35_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_35_lo_lo_hi_lo = {wire_res_70_18,wire_res_70_17,wire_res_70_16,wire_res_70_15,wire_res_70_14,
    wire_res_70_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_35_lo_lo = {wire_res_70_25,wire_res_70_24,wire_res_70_23,wire_res_70_22,wire_res_70_21,
    wire_res_70_20,wire_res_70_19,result_reg_r_35_lo_lo_hi_lo,result_reg_r_35_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_35_lo_hi_lo_lo = {wire_res_70_31,wire_res_70_30,wire_res_70_29,wire_res_70_28,wire_res_70_27,
    wire_res_70_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_35_lo_hi_lo = {wire_res_70_38,wire_res_70_37,wire_res_70_36,wire_res_70_35,wire_res_70_34,
    wire_res_70_33,wire_res_70_32,result_reg_r_35_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_35_lo_hi_hi_lo = {wire_res_70_45,wire_res_70_44,wire_res_70_43,wire_res_70_42,wire_res_70_41,
    wire_res_70_40,wire_res_70_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_35_lo = {wire_res_70_52,wire_res_70_51,wire_res_70_50,wire_res_70_49,wire_res_70_48,
    wire_res_70_47,wire_res_70_46,result_reg_r_35_lo_hi_hi_lo,result_reg_r_35_lo_hi_lo,result_reg_r_35_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_35_hi_lo_lo_lo = {wire_res_70_58,wire_res_70_57,wire_res_70_56,wire_res_70_55,wire_res_70_54,
    wire_res_70_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_35_hi_lo_lo = {wire_res_70_65,wire_res_70_64,wire_res_70_63,wire_res_70_62,wire_res_70_61,
    wire_res_70_60,wire_res_70_59,result_reg_r_35_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_35_hi_lo_hi_lo = {wire_res_70_71,wire_res_70_70,wire_res_70_69,wire_res_70_68,wire_res_70_67,
    wire_res_70_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_35_hi_lo = {wire_res_70_78,wire_res_70_77,wire_res_70_76,wire_res_70_75,wire_res_70_74,
    wire_res_70_73,wire_res_70_72,result_reg_r_35_hi_lo_hi_lo,result_reg_r_35_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_35_hi_hi_lo_lo = {wire_res_70_84,wire_res_70_83,wire_res_70_82,wire_res_70_81,wire_res_70_80,
    wire_res_70_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_35_hi_hi_lo = {wire_res_70_91,wire_res_70_90,wire_res_70_89,wire_res_70_88,wire_res_70_87,
    wire_res_70_86,wire_res_70_85,result_reg_r_35_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_35_hi_hi_hi_lo = {wire_res_70_98,wire_res_70_97,wire_res_70_96,wire_res_70_95,wire_res_70_94,
    wire_res_70_93,wire_res_70_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_35_hi = {wire_res_70_105,wire_res_70_104,wire_res_70_103,wire_res_70_102,wire_res_70_101,
    wire_res_70_100,wire_res_70_99,result_reg_r_35_hi_hi_hi_lo,result_reg_r_35_hi_hi_lo,result_reg_r_35_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_35_T = {result_reg_r_35_hi,result_reg_r_35_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [138:0] _a_aux_reg_w_36_T_2 = _GEN_1307 - _T_11380; // @[BinaryDesigns2.scala 225:48]
  wire [138:0] _GEN_144 = wire_res_71_33 ? _a_aux_reg_w_36_T_2 : {{33'd0}, a_aux_reg_r_35}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [137:0] _T_11382 = {b_aux_reg_r_35, 32'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_36 = _GEN_144[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [137:0] _GEN_1432 = {{32'd0}, a_aux_reg_w_36}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_72_32 = _GEN_1432 >= _T_11382; // @[BinaryDesigns2.scala 224:35]
  wire [137:0] _a_aux_reg_r_36_T_2 = _GEN_1432 - _T_11382; // @[BinaryDesigns2.scala 225:48]
  wire [137:0] _GEN_146 = wire_res_72_32 ? _a_aux_reg_r_36_T_2 : {{32'd0}, a_aux_reg_w_36}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_36_lo_lo_lo_lo = {wire_res_72_5,wire_res_72_4,wire_res_72_3,wire_res_72_2,wire_res_72_1,
    wire_res_72_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_36_lo_lo_lo = {wire_res_72_12,wire_res_72_11,wire_res_72_10,wire_res_72_9,wire_res_72_8,
    wire_res_72_7,wire_res_72_6,result_reg_r_36_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_36_lo_lo_hi_lo = {wire_res_72_18,wire_res_72_17,wire_res_72_16,wire_res_72_15,wire_res_72_14,
    wire_res_72_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_36_lo_lo = {wire_res_72_25,wire_res_72_24,wire_res_72_23,wire_res_72_22,wire_res_72_21,
    wire_res_72_20,wire_res_72_19,result_reg_r_36_lo_lo_hi_lo,result_reg_r_36_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_36_lo_hi_lo_lo = {wire_res_72_31,wire_res_72_30,wire_res_72_29,wire_res_72_28,wire_res_72_27,
    wire_res_72_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_36_lo_hi_lo = {wire_res_72_38,wire_res_72_37,wire_res_72_36,wire_res_72_35,wire_res_72_34,
    wire_res_72_33,wire_res_72_32,result_reg_r_36_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_36_lo_hi_hi_lo = {wire_res_72_45,wire_res_72_44,wire_res_72_43,wire_res_72_42,wire_res_72_41,
    wire_res_72_40,wire_res_72_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_36_lo = {wire_res_72_52,wire_res_72_51,wire_res_72_50,wire_res_72_49,wire_res_72_48,
    wire_res_72_47,wire_res_72_46,result_reg_r_36_lo_hi_hi_lo,result_reg_r_36_lo_hi_lo,result_reg_r_36_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_36_hi_lo_lo_lo = {wire_res_72_58,wire_res_72_57,wire_res_72_56,wire_res_72_55,wire_res_72_54,
    wire_res_72_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_36_hi_lo_lo = {wire_res_72_65,wire_res_72_64,wire_res_72_63,wire_res_72_62,wire_res_72_61,
    wire_res_72_60,wire_res_72_59,result_reg_r_36_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_36_hi_lo_hi_lo = {wire_res_72_71,wire_res_72_70,wire_res_72_69,wire_res_72_68,wire_res_72_67,
    wire_res_72_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_36_hi_lo = {wire_res_72_78,wire_res_72_77,wire_res_72_76,wire_res_72_75,wire_res_72_74,
    wire_res_72_73,wire_res_72_72,result_reg_r_36_hi_lo_hi_lo,result_reg_r_36_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_36_hi_hi_lo_lo = {wire_res_72_84,wire_res_72_83,wire_res_72_82,wire_res_72_81,wire_res_72_80,
    wire_res_72_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_36_hi_hi_lo = {wire_res_72_91,wire_res_72_90,wire_res_72_89,wire_res_72_88,wire_res_72_87,
    wire_res_72_86,wire_res_72_85,result_reg_r_36_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_36_hi_hi_hi_lo = {wire_res_72_98,wire_res_72_97,wire_res_72_96,wire_res_72_95,wire_res_72_94,
    wire_res_72_93,wire_res_72_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_36_hi = {wire_res_72_105,wire_res_72_104,wire_res_72_103,wire_res_72_102,wire_res_72_101,
    wire_res_72_100,wire_res_72_99,result_reg_r_36_hi_hi_hi_lo,result_reg_r_36_hi_hi_lo,result_reg_r_36_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_36_T = {result_reg_r_36_hi,result_reg_r_36_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [136:0] _a_aux_reg_w_37_T_2 = _GEN_1308 - _T_11384; // @[BinaryDesigns2.scala 225:48]
  wire [136:0] _GEN_148 = wire_res_73_31 ? _a_aux_reg_w_37_T_2 : {{31'd0}, a_aux_reg_r_36}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [135:0] _T_11386 = {b_aux_reg_r_36, 30'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_37 = _GEN_148[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [135:0] _GEN_1435 = {{30'd0}, a_aux_reg_w_37}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_74_30 = _GEN_1435 >= _T_11386; // @[BinaryDesigns2.scala 224:35]
  wire [135:0] _a_aux_reg_r_37_T_2 = _GEN_1435 - _T_11386; // @[BinaryDesigns2.scala 225:48]
  wire [135:0] _GEN_150 = wire_res_74_30 ? _a_aux_reg_r_37_T_2 : {{30'd0}, a_aux_reg_w_37}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_37_lo_lo_lo_lo = {wire_res_74_5,wire_res_74_4,wire_res_74_3,wire_res_74_2,wire_res_74_1,
    wire_res_74_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_37_lo_lo_lo = {wire_res_74_12,wire_res_74_11,wire_res_74_10,wire_res_74_9,wire_res_74_8,
    wire_res_74_7,wire_res_74_6,result_reg_r_37_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_37_lo_lo_hi_lo = {wire_res_74_18,wire_res_74_17,wire_res_74_16,wire_res_74_15,wire_res_74_14,
    wire_res_74_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_37_lo_lo = {wire_res_74_25,wire_res_74_24,wire_res_74_23,wire_res_74_22,wire_res_74_21,
    wire_res_74_20,wire_res_74_19,result_reg_r_37_lo_lo_hi_lo,result_reg_r_37_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_37_lo_hi_lo_lo = {wire_res_74_31,wire_res_74_30,wire_res_74_29,wire_res_74_28,wire_res_74_27,
    wire_res_74_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_37_lo_hi_lo = {wire_res_74_38,wire_res_74_37,wire_res_74_36,wire_res_74_35,wire_res_74_34,
    wire_res_74_33,wire_res_74_32,result_reg_r_37_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_37_lo_hi_hi_lo = {wire_res_74_45,wire_res_74_44,wire_res_74_43,wire_res_74_42,wire_res_74_41,
    wire_res_74_40,wire_res_74_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_37_lo = {wire_res_74_52,wire_res_74_51,wire_res_74_50,wire_res_74_49,wire_res_74_48,
    wire_res_74_47,wire_res_74_46,result_reg_r_37_lo_hi_hi_lo,result_reg_r_37_lo_hi_lo,result_reg_r_37_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_37_hi_lo_lo_lo = {wire_res_74_58,wire_res_74_57,wire_res_74_56,wire_res_74_55,wire_res_74_54,
    wire_res_74_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_37_hi_lo_lo = {wire_res_74_65,wire_res_74_64,wire_res_74_63,wire_res_74_62,wire_res_74_61,
    wire_res_74_60,wire_res_74_59,result_reg_r_37_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_37_hi_lo_hi_lo = {wire_res_74_71,wire_res_74_70,wire_res_74_69,wire_res_74_68,wire_res_74_67,
    wire_res_74_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_37_hi_lo = {wire_res_74_78,wire_res_74_77,wire_res_74_76,wire_res_74_75,wire_res_74_74,
    wire_res_74_73,wire_res_74_72,result_reg_r_37_hi_lo_hi_lo,result_reg_r_37_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_37_hi_hi_lo_lo = {wire_res_74_84,wire_res_74_83,wire_res_74_82,wire_res_74_81,wire_res_74_80,
    wire_res_74_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_37_hi_hi_lo = {wire_res_74_91,wire_res_74_90,wire_res_74_89,wire_res_74_88,wire_res_74_87,
    wire_res_74_86,wire_res_74_85,result_reg_r_37_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_37_hi_hi_hi_lo = {wire_res_74_98,wire_res_74_97,wire_res_74_96,wire_res_74_95,wire_res_74_94,
    wire_res_74_93,wire_res_74_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_37_hi = {wire_res_74_105,wire_res_74_104,wire_res_74_103,wire_res_74_102,wire_res_74_101,
    wire_res_74_100,wire_res_74_99,result_reg_r_37_hi_hi_hi_lo,result_reg_r_37_hi_hi_lo,result_reg_r_37_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_37_T = {result_reg_r_37_hi,result_reg_r_37_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [134:0] _a_aux_reg_w_38_T_2 = _GEN_1309 - _T_11388; // @[BinaryDesigns2.scala 225:48]
  wire [134:0] _GEN_152 = wire_res_75_29 ? _a_aux_reg_w_38_T_2 : {{29'd0}, a_aux_reg_r_37}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [133:0] _T_11390 = {b_aux_reg_r_37, 28'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_38 = _GEN_152[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [133:0] _GEN_1438 = {{28'd0}, a_aux_reg_w_38}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_76_28 = _GEN_1438 >= _T_11390; // @[BinaryDesigns2.scala 224:35]
  wire [133:0] _a_aux_reg_r_38_T_2 = _GEN_1438 - _T_11390; // @[BinaryDesigns2.scala 225:48]
  wire [133:0] _GEN_154 = wire_res_76_28 ? _a_aux_reg_r_38_T_2 : {{28'd0}, a_aux_reg_w_38}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_38_lo_lo_lo_lo = {wire_res_76_5,wire_res_76_4,wire_res_76_3,wire_res_76_2,wire_res_76_1,
    wire_res_76_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_38_lo_lo_lo = {wire_res_76_12,wire_res_76_11,wire_res_76_10,wire_res_76_9,wire_res_76_8,
    wire_res_76_7,wire_res_76_6,result_reg_r_38_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_38_lo_lo_hi_lo = {wire_res_76_18,wire_res_76_17,wire_res_76_16,wire_res_76_15,wire_res_76_14,
    wire_res_76_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_38_lo_lo = {wire_res_76_25,wire_res_76_24,wire_res_76_23,wire_res_76_22,wire_res_76_21,
    wire_res_76_20,wire_res_76_19,result_reg_r_38_lo_lo_hi_lo,result_reg_r_38_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_38_lo_hi_lo_lo = {wire_res_76_31,wire_res_76_30,wire_res_76_29,wire_res_76_28,wire_res_76_27,
    wire_res_76_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_38_lo_hi_lo = {wire_res_76_38,wire_res_76_37,wire_res_76_36,wire_res_76_35,wire_res_76_34,
    wire_res_76_33,wire_res_76_32,result_reg_r_38_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_38_lo_hi_hi_lo = {wire_res_76_45,wire_res_76_44,wire_res_76_43,wire_res_76_42,wire_res_76_41,
    wire_res_76_40,wire_res_76_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_38_lo = {wire_res_76_52,wire_res_76_51,wire_res_76_50,wire_res_76_49,wire_res_76_48,
    wire_res_76_47,wire_res_76_46,result_reg_r_38_lo_hi_hi_lo,result_reg_r_38_lo_hi_lo,result_reg_r_38_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_38_hi_lo_lo_lo = {wire_res_76_58,wire_res_76_57,wire_res_76_56,wire_res_76_55,wire_res_76_54,
    wire_res_76_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_38_hi_lo_lo = {wire_res_76_65,wire_res_76_64,wire_res_76_63,wire_res_76_62,wire_res_76_61,
    wire_res_76_60,wire_res_76_59,result_reg_r_38_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_38_hi_lo_hi_lo = {wire_res_76_71,wire_res_76_70,wire_res_76_69,wire_res_76_68,wire_res_76_67,
    wire_res_76_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_38_hi_lo = {wire_res_76_78,wire_res_76_77,wire_res_76_76,wire_res_76_75,wire_res_76_74,
    wire_res_76_73,wire_res_76_72,result_reg_r_38_hi_lo_hi_lo,result_reg_r_38_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_38_hi_hi_lo_lo = {wire_res_76_84,wire_res_76_83,wire_res_76_82,wire_res_76_81,wire_res_76_80,
    wire_res_76_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_38_hi_hi_lo = {wire_res_76_91,wire_res_76_90,wire_res_76_89,wire_res_76_88,wire_res_76_87,
    wire_res_76_86,wire_res_76_85,result_reg_r_38_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_38_hi_hi_hi_lo = {wire_res_76_98,wire_res_76_97,wire_res_76_96,wire_res_76_95,wire_res_76_94,
    wire_res_76_93,wire_res_76_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_38_hi = {wire_res_76_105,wire_res_76_104,wire_res_76_103,wire_res_76_102,wire_res_76_101,
    wire_res_76_100,wire_res_76_99,result_reg_r_38_hi_hi_hi_lo,result_reg_r_38_hi_hi_lo,result_reg_r_38_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_38_T = {result_reg_r_38_hi,result_reg_r_38_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [132:0] _a_aux_reg_w_39_T_2 = _GEN_1310 - _T_11392; // @[BinaryDesigns2.scala 225:48]
  wire [132:0] _GEN_156 = wire_res_77_27 ? _a_aux_reg_w_39_T_2 : {{27'd0}, a_aux_reg_r_38}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [131:0] _T_11394 = {b_aux_reg_r_38, 26'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_39 = _GEN_156[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [131:0] _GEN_1441 = {{26'd0}, a_aux_reg_w_39}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_78_26 = _GEN_1441 >= _T_11394; // @[BinaryDesigns2.scala 224:35]
  wire [131:0] _a_aux_reg_r_39_T_2 = _GEN_1441 - _T_11394; // @[BinaryDesigns2.scala 225:48]
  wire [131:0] _GEN_158 = wire_res_78_26 ? _a_aux_reg_r_39_T_2 : {{26'd0}, a_aux_reg_w_39}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_39_lo_lo_lo_lo = {wire_res_78_5,wire_res_78_4,wire_res_78_3,wire_res_78_2,wire_res_78_1,
    wire_res_78_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_39_lo_lo_lo = {wire_res_78_12,wire_res_78_11,wire_res_78_10,wire_res_78_9,wire_res_78_8,
    wire_res_78_7,wire_res_78_6,result_reg_r_39_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_39_lo_lo_hi_lo = {wire_res_78_18,wire_res_78_17,wire_res_78_16,wire_res_78_15,wire_res_78_14,
    wire_res_78_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_39_lo_lo = {wire_res_78_25,wire_res_78_24,wire_res_78_23,wire_res_78_22,wire_res_78_21,
    wire_res_78_20,wire_res_78_19,result_reg_r_39_lo_lo_hi_lo,result_reg_r_39_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_39_lo_hi_lo_lo = {wire_res_78_31,wire_res_78_30,wire_res_78_29,wire_res_78_28,wire_res_78_27,
    wire_res_78_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_39_lo_hi_lo = {wire_res_78_38,wire_res_78_37,wire_res_78_36,wire_res_78_35,wire_res_78_34,
    wire_res_78_33,wire_res_78_32,result_reg_r_39_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_39_lo_hi_hi_lo = {wire_res_78_45,wire_res_78_44,wire_res_78_43,wire_res_78_42,wire_res_78_41,
    wire_res_78_40,wire_res_78_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_39_lo = {wire_res_78_52,wire_res_78_51,wire_res_78_50,wire_res_78_49,wire_res_78_48,
    wire_res_78_47,wire_res_78_46,result_reg_r_39_lo_hi_hi_lo,result_reg_r_39_lo_hi_lo,result_reg_r_39_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_39_hi_lo_lo_lo = {wire_res_78_58,wire_res_78_57,wire_res_78_56,wire_res_78_55,wire_res_78_54,
    wire_res_78_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_39_hi_lo_lo = {wire_res_78_65,wire_res_78_64,wire_res_78_63,wire_res_78_62,wire_res_78_61,
    wire_res_78_60,wire_res_78_59,result_reg_r_39_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_39_hi_lo_hi_lo = {wire_res_78_71,wire_res_78_70,wire_res_78_69,wire_res_78_68,wire_res_78_67,
    wire_res_78_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_39_hi_lo = {wire_res_78_78,wire_res_78_77,wire_res_78_76,wire_res_78_75,wire_res_78_74,
    wire_res_78_73,wire_res_78_72,result_reg_r_39_hi_lo_hi_lo,result_reg_r_39_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_39_hi_hi_lo_lo = {wire_res_78_84,wire_res_78_83,wire_res_78_82,wire_res_78_81,wire_res_78_80,
    wire_res_78_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_39_hi_hi_lo = {wire_res_78_91,wire_res_78_90,wire_res_78_89,wire_res_78_88,wire_res_78_87,
    wire_res_78_86,wire_res_78_85,result_reg_r_39_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_39_hi_hi_hi_lo = {wire_res_78_98,wire_res_78_97,wire_res_78_96,wire_res_78_95,wire_res_78_94,
    wire_res_78_93,wire_res_78_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_39_hi = {wire_res_78_105,wire_res_78_104,wire_res_78_103,wire_res_78_102,wire_res_78_101,
    wire_res_78_100,wire_res_78_99,result_reg_r_39_hi_hi_hi_lo,result_reg_r_39_hi_hi_lo,result_reg_r_39_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_39_T = {result_reg_r_39_hi,result_reg_r_39_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [130:0] _a_aux_reg_w_40_T_2 = _GEN_1311 - _T_11396; // @[BinaryDesigns2.scala 225:48]
  wire [130:0] _GEN_160 = wire_res_79_25 ? _a_aux_reg_w_40_T_2 : {{25'd0}, a_aux_reg_r_39}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [129:0] _T_11398 = {b_aux_reg_r_39, 24'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_40 = _GEN_160[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [129:0] _GEN_1444 = {{24'd0}, a_aux_reg_w_40}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_80_24 = _GEN_1444 >= _T_11398; // @[BinaryDesigns2.scala 224:35]
  wire [129:0] _a_aux_reg_r_40_T_2 = _GEN_1444 - _T_11398; // @[BinaryDesigns2.scala 225:48]
  wire [129:0] _GEN_162 = wire_res_80_24 ? _a_aux_reg_r_40_T_2 : {{24'd0}, a_aux_reg_w_40}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_40_lo_lo_lo_lo = {wire_res_80_5,wire_res_80_4,wire_res_80_3,wire_res_80_2,wire_res_80_1,
    wire_res_80_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_40_lo_lo_lo = {wire_res_80_12,wire_res_80_11,wire_res_80_10,wire_res_80_9,wire_res_80_8,
    wire_res_80_7,wire_res_80_6,result_reg_r_40_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_40_lo_lo_hi_lo = {wire_res_80_18,wire_res_80_17,wire_res_80_16,wire_res_80_15,wire_res_80_14,
    wire_res_80_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_40_lo_lo = {wire_res_80_25,wire_res_80_24,wire_res_80_23,wire_res_80_22,wire_res_80_21,
    wire_res_80_20,wire_res_80_19,result_reg_r_40_lo_lo_hi_lo,result_reg_r_40_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_40_lo_hi_lo_lo = {wire_res_80_31,wire_res_80_30,wire_res_80_29,wire_res_80_28,wire_res_80_27,
    wire_res_80_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_40_lo_hi_lo = {wire_res_80_38,wire_res_80_37,wire_res_80_36,wire_res_80_35,wire_res_80_34,
    wire_res_80_33,wire_res_80_32,result_reg_r_40_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_40_lo_hi_hi_lo = {wire_res_80_45,wire_res_80_44,wire_res_80_43,wire_res_80_42,wire_res_80_41,
    wire_res_80_40,wire_res_80_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_40_lo = {wire_res_80_52,wire_res_80_51,wire_res_80_50,wire_res_80_49,wire_res_80_48,
    wire_res_80_47,wire_res_80_46,result_reg_r_40_lo_hi_hi_lo,result_reg_r_40_lo_hi_lo,result_reg_r_40_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_40_hi_lo_lo_lo = {wire_res_80_58,wire_res_80_57,wire_res_80_56,wire_res_80_55,wire_res_80_54,
    wire_res_80_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_40_hi_lo_lo = {wire_res_80_65,wire_res_80_64,wire_res_80_63,wire_res_80_62,wire_res_80_61,
    wire_res_80_60,wire_res_80_59,result_reg_r_40_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_40_hi_lo_hi_lo = {wire_res_80_71,wire_res_80_70,wire_res_80_69,wire_res_80_68,wire_res_80_67,
    wire_res_80_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_40_hi_lo = {wire_res_80_78,wire_res_80_77,wire_res_80_76,wire_res_80_75,wire_res_80_74,
    wire_res_80_73,wire_res_80_72,result_reg_r_40_hi_lo_hi_lo,result_reg_r_40_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_40_hi_hi_lo_lo = {wire_res_80_84,wire_res_80_83,wire_res_80_82,wire_res_80_81,wire_res_80_80,
    wire_res_80_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_40_hi_hi_lo = {wire_res_80_91,wire_res_80_90,wire_res_80_89,wire_res_80_88,wire_res_80_87,
    wire_res_80_86,wire_res_80_85,result_reg_r_40_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_40_hi_hi_hi_lo = {wire_res_80_98,wire_res_80_97,wire_res_80_96,wire_res_80_95,wire_res_80_94,
    wire_res_80_93,wire_res_80_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_40_hi = {wire_res_80_105,wire_res_80_104,wire_res_80_103,wire_res_80_102,wire_res_80_101,
    wire_res_80_100,wire_res_80_99,result_reg_r_40_hi_hi_hi_lo,result_reg_r_40_hi_hi_lo,result_reg_r_40_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_40_T = {result_reg_r_40_hi,result_reg_r_40_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [128:0] _a_aux_reg_w_41_T_2 = _GEN_1312 - _T_11400; // @[BinaryDesigns2.scala 225:48]
  wire [128:0] _GEN_164 = wire_res_81_23 ? _a_aux_reg_w_41_T_2 : {{23'd0}, a_aux_reg_r_40}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [127:0] _T_11402 = {b_aux_reg_r_40, 22'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_41 = _GEN_164[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [127:0] _GEN_1447 = {{22'd0}, a_aux_reg_w_41}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_82_22 = _GEN_1447 >= _T_11402; // @[BinaryDesigns2.scala 224:35]
  wire [127:0] _a_aux_reg_r_41_T_2 = _GEN_1447 - _T_11402; // @[BinaryDesigns2.scala 225:48]
  wire [127:0] _GEN_166 = wire_res_82_22 ? _a_aux_reg_r_41_T_2 : {{22'd0}, a_aux_reg_w_41}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_41_lo_lo_lo_lo = {wire_res_82_5,wire_res_82_4,wire_res_82_3,wire_res_82_2,wire_res_82_1,
    wire_res_82_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_41_lo_lo_lo = {wire_res_82_12,wire_res_82_11,wire_res_82_10,wire_res_82_9,wire_res_82_8,
    wire_res_82_7,wire_res_82_6,result_reg_r_41_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_41_lo_lo_hi_lo = {wire_res_82_18,wire_res_82_17,wire_res_82_16,wire_res_82_15,wire_res_82_14,
    wire_res_82_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_41_lo_lo = {wire_res_82_25,wire_res_82_24,wire_res_82_23,wire_res_82_22,wire_res_82_21,
    wire_res_82_20,wire_res_82_19,result_reg_r_41_lo_lo_hi_lo,result_reg_r_41_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_41_lo_hi_lo_lo = {wire_res_82_31,wire_res_82_30,wire_res_82_29,wire_res_82_28,wire_res_82_27,
    wire_res_82_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_41_lo_hi_lo = {wire_res_82_38,wire_res_82_37,wire_res_82_36,wire_res_82_35,wire_res_82_34,
    wire_res_82_33,wire_res_82_32,result_reg_r_41_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_41_lo_hi_hi_lo = {wire_res_82_45,wire_res_82_44,wire_res_82_43,wire_res_82_42,wire_res_82_41,
    wire_res_82_40,wire_res_82_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_41_lo = {wire_res_82_52,wire_res_82_51,wire_res_82_50,wire_res_82_49,wire_res_82_48,
    wire_res_82_47,wire_res_82_46,result_reg_r_41_lo_hi_hi_lo,result_reg_r_41_lo_hi_lo,result_reg_r_41_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_41_hi_lo_lo_lo = {wire_res_82_58,wire_res_82_57,wire_res_82_56,wire_res_82_55,wire_res_82_54,
    wire_res_82_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_41_hi_lo_lo = {wire_res_82_65,wire_res_82_64,wire_res_82_63,wire_res_82_62,wire_res_82_61,
    wire_res_82_60,wire_res_82_59,result_reg_r_41_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_41_hi_lo_hi_lo = {wire_res_82_71,wire_res_82_70,wire_res_82_69,wire_res_82_68,wire_res_82_67,
    wire_res_82_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_41_hi_lo = {wire_res_82_78,wire_res_82_77,wire_res_82_76,wire_res_82_75,wire_res_82_74,
    wire_res_82_73,wire_res_82_72,result_reg_r_41_hi_lo_hi_lo,result_reg_r_41_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_41_hi_hi_lo_lo = {wire_res_82_84,wire_res_82_83,wire_res_82_82,wire_res_82_81,wire_res_82_80,
    wire_res_82_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_41_hi_hi_lo = {wire_res_82_91,wire_res_82_90,wire_res_82_89,wire_res_82_88,wire_res_82_87,
    wire_res_82_86,wire_res_82_85,result_reg_r_41_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_41_hi_hi_hi_lo = {wire_res_82_98,wire_res_82_97,wire_res_82_96,wire_res_82_95,wire_res_82_94,
    wire_res_82_93,wire_res_82_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_41_hi = {wire_res_82_105,wire_res_82_104,wire_res_82_103,wire_res_82_102,wire_res_82_101,
    wire_res_82_100,wire_res_82_99,result_reg_r_41_hi_hi_hi_lo,result_reg_r_41_hi_hi_lo,result_reg_r_41_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_41_T = {result_reg_r_41_hi,result_reg_r_41_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [126:0] _a_aux_reg_w_42_T_2 = _GEN_1313 - _T_11404; // @[BinaryDesigns2.scala 225:48]
  wire [126:0] _GEN_168 = wire_res_83_21 ? _a_aux_reg_w_42_T_2 : {{21'd0}, a_aux_reg_r_41}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [125:0] _T_11406 = {b_aux_reg_r_41, 20'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_42 = _GEN_168[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [125:0] _GEN_1450 = {{20'd0}, a_aux_reg_w_42}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_84_20 = _GEN_1450 >= _T_11406; // @[BinaryDesigns2.scala 224:35]
  wire [125:0] _a_aux_reg_r_42_T_2 = _GEN_1450 - _T_11406; // @[BinaryDesigns2.scala 225:48]
  wire [125:0] _GEN_170 = wire_res_84_20 ? _a_aux_reg_r_42_T_2 : {{20'd0}, a_aux_reg_w_42}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_42_lo_lo_lo_lo = {wire_res_84_5,wire_res_84_4,wire_res_84_3,wire_res_84_2,wire_res_84_1,
    wire_res_84_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_42_lo_lo_lo = {wire_res_84_12,wire_res_84_11,wire_res_84_10,wire_res_84_9,wire_res_84_8,
    wire_res_84_7,wire_res_84_6,result_reg_r_42_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_42_lo_lo_hi_lo = {wire_res_84_18,wire_res_84_17,wire_res_84_16,wire_res_84_15,wire_res_84_14,
    wire_res_84_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_42_lo_lo = {wire_res_84_25,wire_res_84_24,wire_res_84_23,wire_res_84_22,wire_res_84_21,
    wire_res_84_20,wire_res_84_19,result_reg_r_42_lo_lo_hi_lo,result_reg_r_42_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_42_lo_hi_lo_lo = {wire_res_84_31,wire_res_84_30,wire_res_84_29,wire_res_84_28,wire_res_84_27,
    wire_res_84_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_42_lo_hi_lo = {wire_res_84_38,wire_res_84_37,wire_res_84_36,wire_res_84_35,wire_res_84_34,
    wire_res_84_33,wire_res_84_32,result_reg_r_42_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_42_lo_hi_hi_lo = {wire_res_84_45,wire_res_84_44,wire_res_84_43,wire_res_84_42,wire_res_84_41,
    wire_res_84_40,wire_res_84_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_42_lo = {wire_res_84_52,wire_res_84_51,wire_res_84_50,wire_res_84_49,wire_res_84_48,
    wire_res_84_47,wire_res_84_46,result_reg_r_42_lo_hi_hi_lo,result_reg_r_42_lo_hi_lo,result_reg_r_42_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_42_hi_lo_lo_lo = {wire_res_84_58,wire_res_84_57,wire_res_84_56,wire_res_84_55,wire_res_84_54,
    wire_res_84_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_42_hi_lo_lo = {wire_res_84_65,wire_res_84_64,wire_res_84_63,wire_res_84_62,wire_res_84_61,
    wire_res_84_60,wire_res_84_59,result_reg_r_42_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_42_hi_lo_hi_lo = {wire_res_84_71,wire_res_84_70,wire_res_84_69,wire_res_84_68,wire_res_84_67,
    wire_res_84_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_42_hi_lo = {wire_res_84_78,wire_res_84_77,wire_res_84_76,wire_res_84_75,wire_res_84_74,
    wire_res_84_73,wire_res_84_72,result_reg_r_42_hi_lo_hi_lo,result_reg_r_42_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_42_hi_hi_lo_lo = {wire_res_84_84,wire_res_84_83,wire_res_84_82,wire_res_84_81,wire_res_84_80,
    wire_res_84_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_42_hi_hi_lo = {wire_res_84_91,wire_res_84_90,wire_res_84_89,wire_res_84_88,wire_res_84_87,
    wire_res_84_86,wire_res_84_85,result_reg_r_42_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_42_hi_hi_hi_lo = {wire_res_84_98,wire_res_84_97,wire_res_84_96,wire_res_84_95,wire_res_84_94,
    wire_res_84_93,wire_res_84_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_42_hi = {wire_res_84_105,wire_res_84_104,wire_res_84_103,wire_res_84_102,wire_res_84_101,
    wire_res_84_100,wire_res_84_99,result_reg_r_42_hi_hi_hi_lo,result_reg_r_42_hi_hi_lo,result_reg_r_42_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_42_T = {result_reg_r_42_hi,result_reg_r_42_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [124:0] _a_aux_reg_w_43_T_2 = _GEN_1314 - _T_11408; // @[BinaryDesigns2.scala 225:48]
  wire [124:0] _GEN_172 = wire_res_85_19 ? _a_aux_reg_w_43_T_2 : {{19'd0}, a_aux_reg_r_42}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [123:0] _T_11410 = {b_aux_reg_r_42, 18'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_43 = _GEN_172[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [123:0] _GEN_1453 = {{18'd0}, a_aux_reg_w_43}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_86_18 = _GEN_1453 >= _T_11410; // @[BinaryDesigns2.scala 224:35]
  wire [123:0] _a_aux_reg_r_43_T_2 = _GEN_1453 - _T_11410; // @[BinaryDesigns2.scala 225:48]
  wire [123:0] _GEN_174 = wire_res_86_18 ? _a_aux_reg_r_43_T_2 : {{18'd0}, a_aux_reg_w_43}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_43_lo_lo_lo_lo = {wire_res_86_5,wire_res_86_4,wire_res_86_3,wire_res_86_2,wire_res_86_1,
    wire_res_86_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_43_lo_lo_lo = {wire_res_86_12,wire_res_86_11,wire_res_86_10,wire_res_86_9,wire_res_86_8,
    wire_res_86_7,wire_res_86_6,result_reg_r_43_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_43_lo_lo_hi_lo = {wire_res_86_18,wire_res_86_17,wire_res_86_16,wire_res_86_15,wire_res_86_14,
    wire_res_86_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_43_lo_lo = {wire_res_86_25,wire_res_86_24,wire_res_86_23,wire_res_86_22,wire_res_86_21,
    wire_res_86_20,wire_res_86_19,result_reg_r_43_lo_lo_hi_lo,result_reg_r_43_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_43_lo_hi_lo_lo = {wire_res_86_31,wire_res_86_30,wire_res_86_29,wire_res_86_28,wire_res_86_27,
    wire_res_86_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_43_lo_hi_lo = {wire_res_86_38,wire_res_86_37,wire_res_86_36,wire_res_86_35,wire_res_86_34,
    wire_res_86_33,wire_res_86_32,result_reg_r_43_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_43_lo_hi_hi_lo = {wire_res_86_45,wire_res_86_44,wire_res_86_43,wire_res_86_42,wire_res_86_41,
    wire_res_86_40,wire_res_86_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_43_lo = {wire_res_86_52,wire_res_86_51,wire_res_86_50,wire_res_86_49,wire_res_86_48,
    wire_res_86_47,wire_res_86_46,result_reg_r_43_lo_hi_hi_lo,result_reg_r_43_lo_hi_lo,result_reg_r_43_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_43_hi_lo_lo_lo = {wire_res_86_58,wire_res_86_57,wire_res_86_56,wire_res_86_55,wire_res_86_54,
    wire_res_86_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_43_hi_lo_lo = {wire_res_86_65,wire_res_86_64,wire_res_86_63,wire_res_86_62,wire_res_86_61,
    wire_res_86_60,wire_res_86_59,result_reg_r_43_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_43_hi_lo_hi_lo = {wire_res_86_71,wire_res_86_70,wire_res_86_69,wire_res_86_68,wire_res_86_67,
    wire_res_86_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_43_hi_lo = {wire_res_86_78,wire_res_86_77,wire_res_86_76,wire_res_86_75,wire_res_86_74,
    wire_res_86_73,wire_res_86_72,result_reg_r_43_hi_lo_hi_lo,result_reg_r_43_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_43_hi_hi_lo_lo = {wire_res_86_84,wire_res_86_83,wire_res_86_82,wire_res_86_81,wire_res_86_80,
    wire_res_86_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_43_hi_hi_lo = {wire_res_86_91,wire_res_86_90,wire_res_86_89,wire_res_86_88,wire_res_86_87,
    wire_res_86_86,wire_res_86_85,result_reg_r_43_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_43_hi_hi_hi_lo = {wire_res_86_98,wire_res_86_97,wire_res_86_96,wire_res_86_95,wire_res_86_94,
    wire_res_86_93,wire_res_86_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_43_hi = {wire_res_86_105,wire_res_86_104,wire_res_86_103,wire_res_86_102,wire_res_86_101,
    wire_res_86_100,wire_res_86_99,result_reg_r_43_hi_hi_hi_lo,result_reg_r_43_hi_hi_lo,result_reg_r_43_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_43_T = {result_reg_r_43_hi,result_reg_r_43_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [122:0] _a_aux_reg_w_44_T_2 = _GEN_1315 - _T_11412; // @[BinaryDesigns2.scala 225:48]
  wire [122:0] _GEN_176 = wire_res_87_17 ? _a_aux_reg_w_44_T_2 : {{17'd0}, a_aux_reg_r_43}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [121:0] _T_11414 = {b_aux_reg_r_43, 16'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_44 = _GEN_176[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [121:0] _GEN_1456 = {{16'd0}, a_aux_reg_w_44}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_88_16 = _GEN_1456 >= _T_11414; // @[BinaryDesigns2.scala 224:35]
  wire [121:0] _a_aux_reg_r_44_T_2 = _GEN_1456 - _T_11414; // @[BinaryDesigns2.scala 225:48]
  wire [121:0] _GEN_178 = wire_res_88_16 ? _a_aux_reg_r_44_T_2 : {{16'd0}, a_aux_reg_w_44}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_44_lo_lo_lo_lo = {wire_res_88_5,wire_res_88_4,wire_res_88_3,wire_res_88_2,wire_res_88_1,
    wire_res_88_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_44_lo_lo_lo = {wire_res_88_12,wire_res_88_11,wire_res_88_10,wire_res_88_9,wire_res_88_8,
    wire_res_88_7,wire_res_88_6,result_reg_r_44_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_44_lo_lo_hi_lo = {wire_res_88_18,wire_res_88_17,wire_res_88_16,wire_res_88_15,wire_res_88_14,
    wire_res_88_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_44_lo_lo = {wire_res_88_25,wire_res_88_24,wire_res_88_23,wire_res_88_22,wire_res_88_21,
    wire_res_88_20,wire_res_88_19,result_reg_r_44_lo_lo_hi_lo,result_reg_r_44_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_44_lo_hi_lo_lo = {wire_res_88_31,wire_res_88_30,wire_res_88_29,wire_res_88_28,wire_res_88_27,
    wire_res_88_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_44_lo_hi_lo = {wire_res_88_38,wire_res_88_37,wire_res_88_36,wire_res_88_35,wire_res_88_34,
    wire_res_88_33,wire_res_88_32,result_reg_r_44_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_44_lo_hi_hi_lo = {wire_res_88_45,wire_res_88_44,wire_res_88_43,wire_res_88_42,wire_res_88_41,
    wire_res_88_40,wire_res_88_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_44_lo = {wire_res_88_52,wire_res_88_51,wire_res_88_50,wire_res_88_49,wire_res_88_48,
    wire_res_88_47,wire_res_88_46,result_reg_r_44_lo_hi_hi_lo,result_reg_r_44_lo_hi_lo,result_reg_r_44_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_44_hi_lo_lo_lo = {wire_res_88_58,wire_res_88_57,wire_res_88_56,wire_res_88_55,wire_res_88_54,
    wire_res_88_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_44_hi_lo_lo = {wire_res_88_65,wire_res_88_64,wire_res_88_63,wire_res_88_62,wire_res_88_61,
    wire_res_88_60,wire_res_88_59,result_reg_r_44_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_44_hi_lo_hi_lo = {wire_res_88_71,wire_res_88_70,wire_res_88_69,wire_res_88_68,wire_res_88_67,
    wire_res_88_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_44_hi_lo = {wire_res_88_78,wire_res_88_77,wire_res_88_76,wire_res_88_75,wire_res_88_74,
    wire_res_88_73,wire_res_88_72,result_reg_r_44_hi_lo_hi_lo,result_reg_r_44_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_44_hi_hi_lo_lo = {wire_res_88_84,wire_res_88_83,wire_res_88_82,wire_res_88_81,wire_res_88_80,
    wire_res_88_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_44_hi_hi_lo = {wire_res_88_91,wire_res_88_90,wire_res_88_89,wire_res_88_88,wire_res_88_87,
    wire_res_88_86,wire_res_88_85,result_reg_r_44_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_44_hi_hi_hi_lo = {wire_res_88_98,wire_res_88_97,wire_res_88_96,wire_res_88_95,wire_res_88_94,
    wire_res_88_93,wire_res_88_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_44_hi = {wire_res_88_105,wire_res_88_104,wire_res_88_103,wire_res_88_102,wire_res_88_101,
    wire_res_88_100,wire_res_88_99,result_reg_r_44_hi_hi_hi_lo,result_reg_r_44_hi_hi_lo,result_reg_r_44_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_44_T = {result_reg_r_44_hi,result_reg_r_44_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [120:0] _a_aux_reg_w_45_T_2 = _GEN_1316 - _T_11416; // @[BinaryDesigns2.scala 225:48]
  wire [120:0] _GEN_180 = wire_res_89_15 ? _a_aux_reg_w_45_T_2 : {{15'd0}, a_aux_reg_r_44}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [119:0] _T_11418 = {b_aux_reg_r_44, 14'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_45 = _GEN_180[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [119:0] _GEN_1459 = {{14'd0}, a_aux_reg_w_45}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_90_14 = _GEN_1459 >= _T_11418; // @[BinaryDesigns2.scala 224:35]
  wire [119:0] _a_aux_reg_r_45_T_2 = _GEN_1459 - _T_11418; // @[BinaryDesigns2.scala 225:48]
  wire [119:0] _GEN_182 = wire_res_90_14 ? _a_aux_reg_r_45_T_2 : {{14'd0}, a_aux_reg_w_45}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_45_lo_lo_lo_lo = {wire_res_90_5,wire_res_90_4,wire_res_90_3,wire_res_90_2,wire_res_90_1,
    wire_res_90_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_45_lo_lo_lo = {wire_res_90_12,wire_res_90_11,wire_res_90_10,wire_res_90_9,wire_res_90_8,
    wire_res_90_7,wire_res_90_6,result_reg_r_45_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_45_lo_lo_hi_lo = {wire_res_90_18,wire_res_90_17,wire_res_90_16,wire_res_90_15,wire_res_90_14,
    wire_res_90_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_45_lo_lo = {wire_res_90_25,wire_res_90_24,wire_res_90_23,wire_res_90_22,wire_res_90_21,
    wire_res_90_20,wire_res_90_19,result_reg_r_45_lo_lo_hi_lo,result_reg_r_45_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_45_lo_hi_lo_lo = {wire_res_90_31,wire_res_90_30,wire_res_90_29,wire_res_90_28,wire_res_90_27,
    wire_res_90_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_45_lo_hi_lo = {wire_res_90_38,wire_res_90_37,wire_res_90_36,wire_res_90_35,wire_res_90_34,
    wire_res_90_33,wire_res_90_32,result_reg_r_45_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_45_lo_hi_hi_lo = {wire_res_90_45,wire_res_90_44,wire_res_90_43,wire_res_90_42,wire_res_90_41,
    wire_res_90_40,wire_res_90_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_45_lo = {wire_res_90_52,wire_res_90_51,wire_res_90_50,wire_res_90_49,wire_res_90_48,
    wire_res_90_47,wire_res_90_46,result_reg_r_45_lo_hi_hi_lo,result_reg_r_45_lo_hi_lo,result_reg_r_45_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_45_hi_lo_lo_lo = {wire_res_90_58,wire_res_90_57,wire_res_90_56,wire_res_90_55,wire_res_90_54,
    wire_res_90_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_45_hi_lo_lo = {wire_res_90_65,wire_res_90_64,wire_res_90_63,wire_res_90_62,wire_res_90_61,
    wire_res_90_60,wire_res_90_59,result_reg_r_45_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_45_hi_lo_hi_lo = {wire_res_90_71,wire_res_90_70,wire_res_90_69,wire_res_90_68,wire_res_90_67,
    wire_res_90_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_45_hi_lo = {wire_res_90_78,wire_res_90_77,wire_res_90_76,wire_res_90_75,wire_res_90_74,
    wire_res_90_73,wire_res_90_72,result_reg_r_45_hi_lo_hi_lo,result_reg_r_45_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_45_hi_hi_lo_lo = {wire_res_90_84,wire_res_90_83,wire_res_90_82,wire_res_90_81,wire_res_90_80,
    wire_res_90_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_45_hi_hi_lo = {wire_res_90_91,wire_res_90_90,wire_res_90_89,wire_res_90_88,wire_res_90_87,
    wire_res_90_86,wire_res_90_85,result_reg_r_45_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_45_hi_hi_hi_lo = {wire_res_90_98,wire_res_90_97,wire_res_90_96,wire_res_90_95,wire_res_90_94,
    wire_res_90_93,wire_res_90_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_45_hi = {wire_res_90_105,wire_res_90_104,wire_res_90_103,wire_res_90_102,wire_res_90_101,
    wire_res_90_100,wire_res_90_99,result_reg_r_45_hi_hi_hi_lo,result_reg_r_45_hi_hi_lo,result_reg_r_45_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_45_T = {result_reg_r_45_hi,result_reg_r_45_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [118:0] _a_aux_reg_w_46_T_2 = _GEN_1317 - _T_11420; // @[BinaryDesigns2.scala 225:48]
  wire [118:0] _GEN_184 = wire_res_91_13 ? _a_aux_reg_w_46_T_2 : {{13'd0}, a_aux_reg_r_45}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [117:0] _T_11422 = {b_aux_reg_r_45, 12'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_46 = _GEN_184[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [117:0] _GEN_1462 = {{12'd0}, a_aux_reg_w_46}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_92_12 = _GEN_1462 >= _T_11422; // @[BinaryDesigns2.scala 224:35]
  wire [117:0] _a_aux_reg_r_46_T_2 = _GEN_1462 - _T_11422; // @[BinaryDesigns2.scala 225:48]
  wire [117:0] _GEN_186 = wire_res_92_12 ? _a_aux_reg_r_46_T_2 : {{12'd0}, a_aux_reg_w_46}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_46_lo_lo_lo_lo = {wire_res_92_5,wire_res_92_4,wire_res_92_3,wire_res_92_2,wire_res_92_1,
    wire_res_92_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_46_lo_lo_lo = {wire_res_92_12,wire_res_92_11,wire_res_92_10,wire_res_92_9,wire_res_92_8,
    wire_res_92_7,wire_res_92_6,result_reg_r_46_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_46_lo_lo_hi_lo = {wire_res_92_18,wire_res_92_17,wire_res_92_16,wire_res_92_15,wire_res_92_14,
    wire_res_92_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_46_lo_lo = {wire_res_92_25,wire_res_92_24,wire_res_92_23,wire_res_92_22,wire_res_92_21,
    wire_res_92_20,wire_res_92_19,result_reg_r_46_lo_lo_hi_lo,result_reg_r_46_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_46_lo_hi_lo_lo = {wire_res_92_31,wire_res_92_30,wire_res_92_29,wire_res_92_28,wire_res_92_27,
    wire_res_92_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_46_lo_hi_lo = {wire_res_92_38,wire_res_92_37,wire_res_92_36,wire_res_92_35,wire_res_92_34,
    wire_res_92_33,wire_res_92_32,result_reg_r_46_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_46_lo_hi_hi_lo = {wire_res_92_45,wire_res_92_44,wire_res_92_43,wire_res_92_42,wire_res_92_41,
    wire_res_92_40,wire_res_92_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_46_lo = {wire_res_92_52,wire_res_92_51,wire_res_92_50,wire_res_92_49,wire_res_92_48,
    wire_res_92_47,wire_res_92_46,result_reg_r_46_lo_hi_hi_lo,result_reg_r_46_lo_hi_lo,result_reg_r_46_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_46_hi_lo_lo_lo = {wire_res_92_58,wire_res_92_57,wire_res_92_56,wire_res_92_55,wire_res_92_54,
    wire_res_92_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_46_hi_lo_lo = {wire_res_92_65,wire_res_92_64,wire_res_92_63,wire_res_92_62,wire_res_92_61,
    wire_res_92_60,wire_res_92_59,result_reg_r_46_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_46_hi_lo_hi_lo = {wire_res_92_71,wire_res_92_70,wire_res_92_69,wire_res_92_68,wire_res_92_67,
    wire_res_92_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_46_hi_lo = {wire_res_92_78,wire_res_92_77,wire_res_92_76,wire_res_92_75,wire_res_92_74,
    wire_res_92_73,wire_res_92_72,result_reg_r_46_hi_lo_hi_lo,result_reg_r_46_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_46_hi_hi_lo_lo = {wire_res_92_84,wire_res_92_83,wire_res_92_82,wire_res_92_81,wire_res_92_80,
    wire_res_92_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_46_hi_hi_lo = {wire_res_92_91,wire_res_92_90,wire_res_92_89,wire_res_92_88,wire_res_92_87,
    wire_res_92_86,wire_res_92_85,result_reg_r_46_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_46_hi_hi_hi_lo = {wire_res_92_98,wire_res_92_97,wire_res_92_96,wire_res_92_95,wire_res_92_94,
    wire_res_92_93,wire_res_92_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_46_hi = {wire_res_92_105,wire_res_92_104,wire_res_92_103,wire_res_92_102,wire_res_92_101,
    wire_res_92_100,wire_res_92_99,result_reg_r_46_hi_hi_hi_lo,result_reg_r_46_hi_hi_lo,result_reg_r_46_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_46_T = {result_reg_r_46_hi,result_reg_r_46_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [116:0] _a_aux_reg_w_47_T_2 = _GEN_1318 - _T_11424; // @[BinaryDesigns2.scala 225:48]
  wire [116:0] _GEN_188 = wire_res_93_11 ? _a_aux_reg_w_47_T_2 : {{11'd0}, a_aux_reg_r_46}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [115:0] _T_11426 = {b_aux_reg_r_46, 10'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_47 = _GEN_188[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [115:0] _GEN_1465 = {{10'd0}, a_aux_reg_w_47}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_94_10 = _GEN_1465 >= _T_11426; // @[BinaryDesigns2.scala 224:35]
  wire [115:0] _a_aux_reg_r_47_T_2 = _GEN_1465 - _T_11426; // @[BinaryDesigns2.scala 225:48]
  wire [115:0] _GEN_190 = wire_res_94_10 ? _a_aux_reg_r_47_T_2 : {{10'd0}, a_aux_reg_w_47}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_47_lo_lo_lo_lo = {wire_res_94_5,wire_res_94_4,wire_res_94_3,wire_res_94_2,wire_res_94_1,
    wire_res_94_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_47_lo_lo_lo = {wire_res_94_12,wire_res_94_11,wire_res_94_10,wire_res_94_9,wire_res_94_8,
    wire_res_94_7,wire_res_94_6,result_reg_r_47_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_47_lo_lo_hi_lo = {wire_res_94_18,wire_res_94_17,wire_res_94_16,wire_res_94_15,wire_res_94_14,
    wire_res_94_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_47_lo_lo = {wire_res_94_25,wire_res_94_24,wire_res_94_23,wire_res_94_22,wire_res_94_21,
    wire_res_94_20,wire_res_94_19,result_reg_r_47_lo_lo_hi_lo,result_reg_r_47_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_47_lo_hi_lo_lo = {wire_res_94_31,wire_res_94_30,wire_res_94_29,wire_res_94_28,wire_res_94_27,
    wire_res_94_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_47_lo_hi_lo = {wire_res_94_38,wire_res_94_37,wire_res_94_36,wire_res_94_35,wire_res_94_34,
    wire_res_94_33,wire_res_94_32,result_reg_r_47_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_47_lo_hi_hi_lo = {wire_res_94_45,wire_res_94_44,wire_res_94_43,wire_res_94_42,wire_res_94_41,
    wire_res_94_40,wire_res_94_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_47_lo = {wire_res_94_52,wire_res_94_51,wire_res_94_50,wire_res_94_49,wire_res_94_48,
    wire_res_94_47,wire_res_94_46,result_reg_r_47_lo_hi_hi_lo,result_reg_r_47_lo_hi_lo,result_reg_r_47_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_47_hi_lo_lo_lo = {wire_res_94_58,wire_res_94_57,wire_res_94_56,wire_res_94_55,wire_res_94_54,
    wire_res_94_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_47_hi_lo_lo = {wire_res_94_65,wire_res_94_64,wire_res_94_63,wire_res_94_62,wire_res_94_61,
    wire_res_94_60,wire_res_94_59,result_reg_r_47_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_47_hi_lo_hi_lo = {wire_res_94_71,wire_res_94_70,wire_res_94_69,wire_res_94_68,wire_res_94_67,
    wire_res_94_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_47_hi_lo = {wire_res_94_78,wire_res_94_77,wire_res_94_76,wire_res_94_75,wire_res_94_74,
    wire_res_94_73,wire_res_94_72,result_reg_r_47_hi_lo_hi_lo,result_reg_r_47_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_47_hi_hi_lo_lo = {wire_res_94_84,wire_res_94_83,wire_res_94_82,wire_res_94_81,wire_res_94_80,
    wire_res_94_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_47_hi_hi_lo = {wire_res_94_91,wire_res_94_90,wire_res_94_89,wire_res_94_88,wire_res_94_87,
    wire_res_94_86,wire_res_94_85,result_reg_r_47_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_47_hi_hi_hi_lo = {wire_res_94_98,wire_res_94_97,wire_res_94_96,wire_res_94_95,wire_res_94_94,
    wire_res_94_93,wire_res_94_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_47_hi = {wire_res_94_105,wire_res_94_104,wire_res_94_103,wire_res_94_102,wire_res_94_101,
    wire_res_94_100,wire_res_94_99,result_reg_r_47_hi_hi_hi_lo,result_reg_r_47_hi_hi_lo,result_reg_r_47_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_47_T = {result_reg_r_47_hi,result_reg_r_47_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [114:0] _a_aux_reg_w_48_T_2 = _GEN_1319 - _T_11428; // @[BinaryDesigns2.scala 225:48]
  wire [114:0] _GEN_192 = wire_res_95_9 ? _a_aux_reg_w_48_T_2 : {{9'd0}, a_aux_reg_r_47}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [113:0] _T_11430 = {b_aux_reg_r_47, 8'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_48 = _GEN_192[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [113:0] _GEN_1468 = {{8'd0}, a_aux_reg_w_48}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_96_8 = _GEN_1468 >= _T_11430; // @[BinaryDesigns2.scala 224:35]
  wire [113:0] _a_aux_reg_r_48_T_2 = _GEN_1468 - _T_11430; // @[BinaryDesigns2.scala 225:48]
  wire [113:0] _GEN_194 = wire_res_96_8 ? _a_aux_reg_r_48_T_2 : {{8'd0}, a_aux_reg_w_48}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_48_lo_lo_lo_lo = {wire_res_96_5,wire_res_96_4,wire_res_96_3,wire_res_96_2,wire_res_96_1,
    wire_res_96_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_48_lo_lo_lo = {wire_res_96_12,wire_res_96_11,wire_res_96_10,wire_res_96_9,wire_res_96_8,
    wire_res_96_7,wire_res_96_6,result_reg_r_48_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_48_lo_lo_hi_lo = {wire_res_96_18,wire_res_96_17,wire_res_96_16,wire_res_96_15,wire_res_96_14,
    wire_res_96_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_48_lo_lo = {wire_res_96_25,wire_res_96_24,wire_res_96_23,wire_res_96_22,wire_res_96_21,
    wire_res_96_20,wire_res_96_19,result_reg_r_48_lo_lo_hi_lo,result_reg_r_48_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_48_lo_hi_lo_lo = {wire_res_96_31,wire_res_96_30,wire_res_96_29,wire_res_96_28,wire_res_96_27,
    wire_res_96_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_48_lo_hi_lo = {wire_res_96_38,wire_res_96_37,wire_res_96_36,wire_res_96_35,wire_res_96_34,
    wire_res_96_33,wire_res_96_32,result_reg_r_48_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_48_lo_hi_hi_lo = {wire_res_96_45,wire_res_96_44,wire_res_96_43,wire_res_96_42,wire_res_96_41,
    wire_res_96_40,wire_res_96_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_48_lo = {wire_res_96_52,wire_res_96_51,wire_res_96_50,wire_res_96_49,wire_res_96_48,
    wire_res_96_47,wire_res_96_46,result_reg_r_48_lo_hi_hi_lo,result_reg_r_48_lo_hi_lo,result_reg_r_48_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_48_hi_lo_lo_lo = {wire_res_96_58,wire_res_96_57,wire_res_96_56,wire_res_96_55,wire_res_96_54,
    wire_res_96_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_48_hi_lo_lo = {wire_res_96_65,wire_res_96_64,wire_res_96_63,wire_res_96_62,wire_res_96_61,
    wire_res_96_60,wire_res_96_59,result_reg_r_48_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_48_hi_lo_hi_lo = {wire_res_96_71,wire_res_96_70,wire_res_96_69,wire_res_96_68,wire_res_96_67,
    wire_res_96_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_48_hi_lo = {wire_res_96_78,wire_res_96_77,wire_res_96_76,wire_res_96_75,wire_res_96_74,
    wire_res_96_73,wire_res_96_72,result_reg_r_48_hi_lo_hi_lo,result_reg_r_48_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_48_hi_hi_lo_lo = {wire_res_96_84,wire_res_96_83,wire_res_96_82,wire_res_96_81,wire_res_96_80,
    wire_res_96_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_48_hi_hi_lo = {wire_res_96_91,wire_res_96_90,wire_res_96_89,wire_res_96_88,wire_res_96_87,
    wire_res_96_86,wire_res_96_85,result_reg_r_48_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_48_hi_hi_hi_lo = {wire_res_96_98,wire_res_96_97,wire_res_96_96,wire_res_96_95,wire_res_96_94,
    wire_res_96_93,wire_res_96_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_48_hi = {wire_res_96_105,wire_res_96_104,wire_res_96_103,wire_res_96_102,wire_res_96_101,
    wire_res_96_100,wire_res_96_99,result_reg_r_48_hi_hi_hi_lo,result_reg_r_48_hi_hi_lo,result_reg_r_48_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_48_T = {result_reg_r_48_hi,result_reg_r_48_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [112:0] _a_aux_reg_w_49_T_2 = _GEN_1320 - _T_11432; // @[BinaryDesigns2.scala 225:48]
  wire [112:0] _GEN_196 = wire_res_97_7 ? _a_aux_reg_w_49_T_2 : {{7'd0}, a_aux_reg_r_48}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [111:0] _T_11434 = {b_aux_reg_r_48, 6'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_49 = _GEN_196[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [111:0] _GEN_1471 = {{6'd0}, a_aux_reg_w_49}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_98_6 = _GEN_1471 >= _T_11434; // @[BinaryDesigns2.scala 224:35]
  wire [111:0] _a_aux_reg_r_49_T_2 = _GEN_1471 - _T_11434; // @[BinaryDesigns2.scala 225:48]
  wire [111:0] _GEN_198 = wire_res_98_6 ? _a_aux_reg_r_49_T_2 : {{6'd0}, a_aux_reg_w_49}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_49_lo_lo_lo_lo = {wire_res_98_5,wire_res_98_4,wire_res_98_3,wire_res_98_2,wire_res_98_1,
    wire_res_98_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_49_lo_lo_lo = {wire_res_98_12,wire_res_98_11,wire_res_98_10,wire_res_98_9,wire_res_98_8,
    wire_res_98_7,wire_res_98_6,result_reg_r_49_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_49_lo_lo_hi_lo = {wire_res_98_18,wire_res_98_17,wire_res_98_16,wire_res_98_15,wire_res_98_14,
    wire_res_98_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_49_lo_lo = {wire_res_98_25,wire_res_98_24,wire_res_98_23,wire_res_98_22,wire_res_98_21,
    wire_res_98_20,wire_res_98_19,result_reg_r_49_lo_lo_hi_lo,result_reg_r_49_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_49_lo_hi_lo_lo = {wire_res_98_31,wire_res_98_30,wire_res_98_29,wire_res_98_28,wire_res_98_27,
    wire_res_98_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_49_lo_hi_lo = {wire_res_98_38,wire_res_98_37,wire_res_98_36,wire_res_98_35,wire_res_98_34,
    wire_res_98_33,wire_res_98_32,result_reg_r_49_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_49_lo_hi_hi_lo = {wire_res_98_45,wire_res_98_44,wire_res_98_43,wire_res_98_42,wire_res_98_41,
    wire_res_98_40,wire_res_98_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_49_lo = {wire_res_98_52,wire_res_98_51,wire_res_98_50,wire_res_98_49,wire_res_98_48,
    wire_res_98_47,wire_res_98_46,result_reg_r_49_lo_hi_hi_lo,result_reg_r_49_lo_hi_lo,result_reg_r_49_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_49_hi_lo_lo_lo = {wire_res_98_58,wire_res_98_57,wire_res_98_56,wire_res_98_55,wire_res_98_54,
    wire_res_98_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_49_hi_lo_lo = {wire_res_98_65,wire_res_98_64,wire_res_98_63,wire_res_98_62,wire_res_98_61,
    wire_res_98_60,wire_res_98_59,result_reg_r_49_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_49_hi_lo_hi_lo = {wire_res_98_71,wire_res_98_70,wire_res_98_69,wire_res_98_68,wire_res_98_67,
    wire_res_98_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_49_hi_lo = {wire_res_98_78,wire_res_98_77,wire_res_98_76,wire_res_98_75,wire_res_98_74,
    wire_res_98_73,wire_res_98_72,result_reg_r_49_hi_lo_hi_lo,result_reg_r_49_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_49_hi_hi_lo_lo = {wire_res_98_84,wire_res_98_83,wire_res_98_82,wire_res_98_81,wire_res_98_80,
    wire_res_98_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_49_hi_hi_lo = {wire_res_98_91,wire_res_98_90,wire_res_98_89,wire_res_98_88,wire_res_98_87,
    wire_res_98_86,wire_res_98_85,result_reg_r_49_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_49_hi_hi_hi_lo = {wire_res_98_98,wire_res_98_97,wire_res_98_96,wire_res_98_95,wire_res_98_94,
    wire_res_98_93,wire_res_98_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_49_hi = {wire_res_98_105,wire_res_98_104,wire_res_98_103,wire_res_98_102,wire_res_98_101,
    wire_res_98_100,wire_res_98_99,result_reg_r_49_hi_hi_hi_lo,result_reg_r_49_hi_hi_lo,result_reg_r_49_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_49_T = {result_reg_r_49_hi,result_reg_r_49_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [110:0] _a_aux_reg_w_50_T_2 = _GEN_1321 - _T_11436; // @[BinaryDesigns2.scala 225:48]
  wire [110:0] _GEN_200 = wire_res_99_5 ? _a_aux_reg_w_50_T_2 : {{5'd0}, a_aux_reg_r_49}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [109:0] _T_11438 = {b_aux_reg_r_49, 4'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_50 = _GEN_200[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [109:0] _GEN_1474 = {{4'd0}, a_aux_reg_w_50}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_100_4 = _GEN_1474 >= _T_11438; // @[BinaryDesigns2.scala 224:35]
  wire [109:0] _a_aux_reg_r_50_T_2 = _GEN_1474 - _T_11438; // @[BinaryDesigns2.scala 225:48]
  wire [109:0] _GEN_202 = wire_res_100_4 ? _a_aux_reg_r_50_T_2 : {{4'd0}, a_aux_reg_w_50}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_50_lo_lo_lo_lo = {wire_res_100_5,wire_res_100_4,wire_res_100_3,wire_res_100_2,wire_res_100_1,
    wire_res_100_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_50_lo_lo_lo = {wire_res_100_12,wire_res_100_11,wire_res_100_10,wire_res_100_9,wire_res_100_8,
    wire_res_100_7,wire_res_100_6,result_reg_r_50_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_50_lo_lo_hi_lo = {wire_res_100_18,wire_res_100_17,wire_res_100_16,wire_res_100_15,
    wire_res_100_14,wire_res_100_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_50_lo_lo = {wire_res_100_25,wire_res_100_24,wire_res_100_23,wire_res_100_22,wire_res_100_21,
    wire_res_100_20,wire_res_100_19,result_reg_r_50_lo_lo_hi_lo,result_reg_r_50_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_50_lo_hi_lo_lo = {wire_res_100_31,wire_res_100_30,wire_res_100_29,wire_res_100_28,
    wire_res_100_27,wire_res_100_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_50_lo_hi_lo = {wire_res_100_38,wire_res_100_37,wire_res_100_36,wire_res_100_35,
    wire_res_100_34,wire_res_100_33,wire_res_100_32,result_reg_r_50_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_50_lo_hi_hi_lo = {wire_res_100_45,wire_res_100_44,wire_res_100_43,wire_res_100_42,
    wire_res_100_41,wire_res_100_40,wire_res_100_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_50_lo = {wire_res_100_52,wire_res_100_51,wire_res_100_50,wire_res_100_49,wire_res_100_48,
    wire_res_100_47,wire_res_100_46,result_reg_r_50_lo_hi_hi_lo,result_reg_r_50_lo_hi_lo,result_reg_r_50_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_50_hi_lo_lo_lo = {wire_res_100_58,wire_res_100_57,wire_res_100_56,wire_res_100_55,
    wire_res_100_54,wire_res_100_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_50_hi_lo_lo = {wire_res_100_65,wire_res_100_64,wire_res_100_63,wire_res_100_62,
    wire_res_100_61,wire_res_100_60,wire_res_100_59,result_reg_r_50_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_50_hi_lo_hi_lo = {wire_res_100_71,wire_res_100_70,wire_res_100_69,wire_res_100_68,
    wire_res_100_67,wire_res_100_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_50_hi_lo = {wire_res_100_78,wire_res_100_77,wire_res_100_76,wire_res_100_75,wire_res_100_74,
    wire_res_100_73,wire_res_100_72,result_reg_r_50_hi_lo_hi_lo,result_reg_r_50_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_50_hi_hi_lo_lo = {wire_res_100_84,wire_res_100_83,wire_res_100_82,wire_res_100_81,
    wire_res_100_80,wire_res_100_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_50_hi_hi_lo = {wire_res_100_91,wire_res_100_90,wire_res_100_89,wire_res_100_88,
    wire_res_100_87,wire_res_100_86,wire_res_100_85,result_reg_r_50_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_50_hi_hi_hi_lo = {wire_res_100_98,wire_res_100_97,wire_res_100_96,wire_res_100_95,
    wire_res_100_94,wire_res_100_93,wire_res_100_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_50_hi = {wire_res_100_105,wire_res_100_104,wire_res_100_103,wire_res_100_102,wire_res_100_101
    ,wire_res_100_100,wire_res_100_99,result_reg_r_50_hi_hi_hi_lo,result_reg_r_50_hi_hi_lo,result_reg_r_50_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_50_T = {result_reg_r_50_hi,result_reg_r_50_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [108:0] _a_aux_reg_w_51_T_2 = _GEN_1322 - _T_11440; // @[BinaryDesigns2.scala 225:48]
  wire [108:0] _GEN_204 = wire_res_101_3 ? _a_aux_reg_w_51_T_2 : {{3'd0}, a_aux_reg_r_50}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [107:0] _T_11442 = {b_aux_reg_r_50, 2'h0}; // @[BinaryDesigns2.scala 224:56]
  wire [105:0] a_aux_reg_w_51 = _GEN_204[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire [107:0] _GEN_1477 = {{2'd0}, a_aux_reg_w_51}; // @[BinaryDesigns2.scala 224:35]
  wire  wire_res_102_2 = _GEN_1477 >= _T_11442; // @[BinaryDesigns2.scala 224:35]
  wire [107:0] _a_aux_reg_r_51_T_2 = _GEN_1477 - _T_11442; // @[BinaryDesigns2.scala 225:48]
  wire [107:0] _GEN_206 = wire_res_102_2 ? _a_aux_reg_r_51_T_2 : {{2'd0}, a_aux_reg_w_51}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [5:0] result_reg_r_51_lo_lo_lo_lo = {wire_res_102_5,wire_res_102_4,wire_res_102_3,wire_res_102_2,wire_res_102_1,
    wire_res_102_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_51_lo_lo_lo = {wire_res_102_12,wire_res_102_11,wire_res_102_10,wire_res_102_9,wire_res_102_8,
    wire_res_102_7,wire_res_102_6,result_reg_r_51_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_51_lo_lo_hi_lo = {wire_res_102_18,wire_res_102_17,wire_res_102_16,wire_res_102_15,
    wire_res_102_14,wire_res_102_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_51_lo_lo = {wire_res_102_25,wire_res_102_24,wire_res_102_23,wire_res_102_22,wire_res_102_21,
    wire_res_102_20,wire_res_102_19,result_reg_r_51_lo_lo_hi_lo,result_reg_r_51_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_51_lo_hi_lo_lo = {wire_res_102_31,wire_res_102_30,wire_res_102_29,wire_res_102_28,
    wire_res_102_27,wire_res_102_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_51_lo_hi_lo = {wire_res_102_38,wire_res_102_37,wire_res_102_36,wire_res_102_35,
    wire_res_102_34,wire_res_102_33,wire_res_102_32,result_reg_r_51_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_51_lo_hi_hi_lo = {wire_res_102_45,wire_res_102_44,wire_res_102_43,wire_res_102_42,
    wire_res_102_41,wire_res_102_40,wire_res_102_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_51_lo = {wire_res_102_52,wire_res_102_51,wire_res_102_50,wire_res_102_49,wire_res_102_48,
    wire_res_102_47,wire_res_102_46,result_reg_r_51_lo_hi_hi_lo,result_reg_r_51_lo_hi_lo,result_reg_r_51_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_51_hi_lo_lo_lo = {wire_res_102_58,wire_res_102_57,wire_res_102_56,wire_res_102_55,
    wire_res_102_54,wire_res_102_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_51_hi_lo_lo = {wire_res_102_65,wire_res_102_64,wire_res_102_63,wire_res_102_62,
    wire_res_102_61,wire_res_102_60,wire_res_102_59,result_reg_r_51_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_51_hi_lo_hi_lo = {wire_res_102_71,wire_res_102_70,wire_res_102_69,wire_res_102_68,
    wire_res_102_67,wire_res_102_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_51_hi_lo = {wire_res_102_78,wire_res_102_77,wire_res_102_76,wire_res_102_75,wire_res_102_74,
    wire_res_102_73,wire_res_102_72,result_reg_r_51_hi_lo_hi_lo,result_reg_r_51_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_51_hi_hi_lo_lo = {wire_res_102_84,wire_res_102_83,wire_res_102_82,wire_res_102_81,
    wire_res_102_80,wire_res_102_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_51_hi_hi_lo = {wire_res_102_91,wire_res_102_90,wire_res_102_89,wire_res_102_88,
    wire_res_102_87,wire_res_102_86,wire_res_102_85,result_reg_r_51_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_51_hi_hi_hi_lo = {wire_res_102_98,wire_res_102_97,wire_res_102_96,wire_res_102_95,
    wire_res_102_94,wire_res_102_93,wire_res_102_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_51_hi = {wire_res_102_105,wire_res_102_104,wire_res_102_103,wire_res_102_102,wire_res_102_101
    ,wire_res_102_100,wire_res_102_99,result_reg_r_51_hi_hi_hi_lo,result_reg_r_51_hi_hi_lo,result_reg_r_51_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_51_T = {result_reg_r_51_hi,result_reg_r_51_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [106:0] _a_aux_reg_w_52_T_2 = _GEN_1323 - _T_11444; // @[BinaryDesigns2.scala 225:48]
  wire [106:0] _GEN_208 = wire_res_103_1 ? _a_aux_reg_w_52_T_2 : {{1'd0}, a_aux_reg_r_51}; // @[BinaryDesigns2.scala 224:81 225:28 228:28]
  wire [105:0] a_aux_reg_w_52 = _GEN_208[105:0]; // @[BinaryDesigns2.scala 169:27]
  wire  wire_res_104_0 = a_aux_reg_w_52 >= b_aux_reg_r_51; // @[BinaryDesigns2.scala 224:35]
  wire [5:0] result_reg_r_52_lo_lo_lo_lo = {wire_res_104_5,wire_res_104_4,wire_res_104_3,wire_res_104_2,wire_res_104_1,
    wire_res_104_0}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_52_lo_lo_lo = {wire_res_104_12,wire_res_104_11,wire_res_104_10,wire_res_104_9,wire_res_104_8,
    wire_res_104_7,wire_res_104_6,result_reg_r_52_lo_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_52_lo_lo_hi_lo = {wire_res_104_18,wire_res_104_17,wire_res_104_16,wire_res_104_15,
    wire_res_104_14,wire_res_104_13}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_52_lo_lo = {wire_res_104_25,wire_res_104_24,wire_res_104_23,wire_res_104_22,wire_res_104_21,
    wire_res_104_20,wire_res_104_19,result_reg_r_52_lo_lo_hi_lo,result_reg_r_52_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_52_lo_hi_lo_lo = {wire_res_104_31,wire_res_104_30,wire_res_104_29,wire_res_104_28,
    wire_res_104_27,wire_res_104_26}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_52_lo_hi_lo = {wire_res_104_38,wire_res_104_37,wire_res_104_36,wire_res_104_35,
    wire_res_104_34,wire_res_104_33,wire_res_104_32,result_reg_r_52_lo_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_52_lo_hi_hi_lo = {wire_res_104_45,wire_res_104_44,wire_res_104_43,wire_res_104_42,
    wire_res_104_41,wire_res_104_40,wire_res_104_39}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_52_lo = {wire_res_104_52,wire_res_104_51,wire_res_104_50,wire_res_104_49,wire_res_104_48,
    wire_res_104_47,wire_res_104_46,result_reg_r_52_lo_hi_hi_lo,result_reg_r_52_lo_hi_lo,result_reg_r_52_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_52_hi_lo_lo_lo = {wire_res_104_58,wire_res_104_57,wire_res_104_56,wire_res_104_55,
    wire_res_104_54,wire_res_104_53}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_52_hi_lo_lo = {wire_res_104_65,wire_res_104_64,wire_res_104_63,wire_res_104_62,
    wire_res_104_61,wire_res_104_60,wire_res_104_59,result_reg_r_52_hi_lo_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_52_hi_lo_hi_lo = {wire_res_104_71,wire_res_104_70,wire_res_104_69,wire_res_104_68,
    wire_res_104_67,wire_res_104_66}; // @[BinaryDesigns2.scala 231:46]
  wire [25:0] result_reg_r_52_hi_lo = {wire_res_104_78,wire_res_104_77,wire_res_104_76,wire_res_104_75,wire_res_104_74,
    wire_res_104_73,wire_res_104_72,result_reg_r_52_hi_lo_hi_lo,result_reg_r_52_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [5:0] result_reg_r_52_hi_hi_lo_lo = {wire_res_104_84,wire_res_104_83,wire_res_104_82,wire_res_104_81,
    wire_res_104_80,wire_res_104_79}; // @[BinaryDesigns2.scala 231:46]
  wire [12:0] result_reg_r_52_hi_hi_lo = {wire_res_104_91,wire_res_104_90,wire_res_104_89,wire_res_104_88,
    wire_res_104_87,wire_res_104_86,wire_res_104_85,result_reg_r_52_hi_hi_lo_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [6:0] result_reg_r_52_hi_hi_hi_lo = {wire_res_104_98,wire_res_104_97,wire_res_104_96,wire_res_104_95,
    wire_res_104_94,wire_res_104_93,wire_res_104_92}; // @[BinaryDesigns2.scala 231:46]
  wire [52:0] result_reg_r_52_hi = {wire_res_104_105,wire_res_104_104,wire_res_104_103,wire_res_104_102,wire_res_104_101
    ,wire_res_104_100,wire_res_104_99,result_reg_r_52_hi_hi_hi_lo,result_reg_r_52_hi_hi_lo,result_reg_r_52_hi_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [105:0] _result_reg_r_52_T = {result_reg_r_52_hi,result_reg_r_52_lo}; // @[BinaryDesigns2.scala 231:46]
  wire [209:0] _GEN_1480 = reset ? 210'h0 : _GEN_1325; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [207:0] _GEN_1481 = reset ? 208'h0 : _GEN_6; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [205:0] _GEN_1482 = reset ? 206'h0 : _GEN_10; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [203:0] _GEN_1483 = reset ? 204'h0 : _GEN_14; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [201:0] _GEN_1484 = reset ? 202'h0 : _GEN_18; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [199:0] _GEN_1485 = reset ? 200'h0 : _GEN_22; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [197:0] _GEN_1486 = reset ? 198'h0 : _GEN_26; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [195:0] _GEN_1487 = reset ? 196'h0 : _GEN_30; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [193:0] _GEN_1488 = reset ? 194'h0 : _GEN_34; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [191:0] _GEN_1489 = reset ? 192'h0 : _GEN_38; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [189:0] _GEN_1490 = reset ? 190'h0 : _GEN_42; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [187:0] _GEN_1491 = reset ? 188'h0 : _GEN_46; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [185:0] _GEN_1492 = reset ? 186'h0 : _GEN_50; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [183:0] _GEN_1493 = reset ? 184'h0 : _GEN_54; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [181:0] _GEN_1494 = reset ? 182'h0 : _GEN_58; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [179:0] _GEN_1495 = reset ? 180'h0 : _GEN_62; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [177:0] _GEN_1496 = reset ? 178'h0 : _GEN_66; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [175:0] _GEN_1497 = reset ? 176'h0 : _GEN_70; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [173:0] _GEN_1498 = reset ? 174'h0 : _GEN_74; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [171:0] _GEN_1499 = reset ? 172'h0 : _GEN_78; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [169:0] _GEN_1500 = reset ? 170'h0 : _GEN_82; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [167:0] _GEN_1501 = reset ? 168'h0 : _GEN_86; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [165:0] _GEN_1502 = reset ? 166'h0 : _GEN_90; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [163:0] _GEN_1503 = reset ? 164'h0 : _GEN_94; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [161:0] _GEN_1504 = reset ? 162'h0 : _GEN_98; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [159:0] _GEN_1505 = reset ? 160'h0 : _GEN_102; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [157:0] _GEN_1506 = reset ? 158'h0 : _GEN_106; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [155:0] _GEN_1507 = reset ? 156'h0 : _GEN_110; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [153:0] _GEN_1508 = reset ? 154'h0 : _GEN_114; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [151:0] _GEN_1509 = reset ? 152'h0 : _GEN_118; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [149:0] _GEN_1510 = reset ? 150'h0 : _GEN_122; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [147:0] _GEN_1511 = reset ? 148'h0 : _GEN_126; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [145:0] _GEN_1512 = reset ? 146'h0 : _GEN_130; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [143:0] _GEN_1513 = reset ? 144'h0 : _GEN_134; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [141:0] _GEN_1514 = reset ? 142'h0 : _GEN_138; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [139:0] _GEN_1515 = reset ? 140'h0 : _GEN_142; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [137:0] _GEN_1516 = reset ? 138'h0 : _GEN_146; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [135:0] _GEN_1517 = reset ? 136'h0 : _GEN_150; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [133:0] _GEN_1518 = reset ? 134'h0 : _GEN_154; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [131:0] _GEN_1519 = reset ? 132'h0 : _GEN_158; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [129:0] _GEN_1520 = reset ? 130'h0 : _GEN_162; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [127:0] _GEN_1521 = reset ? 128'h0 : _GEN_166; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [125:0] _GEN_1522 = reset ? 126'h0 : _GEN_170; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [123:0] _GEN_1523 = reset ? 124'h0 : _GEN_174; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [121:0] _GEN_1524 = reset ? 122'h0 : _GEN_178; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [119:0] _GEN_1525 = reset ? 120'h0 : _GEN_182; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [117:0] _GEN_1526 = reset ? 118'h0 : _GEN_186; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [115:0] _GEN_1527 = reset ? 116'h0 : _GEN_190; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [113:0] _GEN_1528 = reset ? 114'h0 : _GEN_194; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [111:0] _GEN_1529 = reset ? 112'h0 : _GEN_198; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [109:0] _GEN_1530 = reset ? 110'h0 : _GEN_202; // @[BinaryDesigns2.scala 171:{30,30}]
  wire [107:0] _GEN_1531 = reset ? 108'h0 : _GEN_206; // @[BinaryDesigns2.scala 171:{30,30}]
  assign io_out_s = result_reg_r_52; // @[BinaryDesigns2.scala 195:14]
  always @(posedge clock) begin
    a_aux_reg_r_0 <= _GEN_1480[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_1 <= _GEN_1481[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_2 <= _GEN_1482[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_3 <= _GEN_1483[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_4 <= _GEN_1484[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_5 <= _GEN_1485[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_6 <= _GEN_1486[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_7 <= _GEN_1487[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_8 <= _GEN_1488[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_9 <= _GEN_1489[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_10 <= _GEN_1490[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_11 <= _GEN_1491[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_12 <= _GEN_1492[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_13 <= _GEN_1493[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_14 <= _GEN_1494[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_15 <= _GEN_1495[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_16 <= _GEN_1496[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_17 <= _GEN_1497[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_18 <= _GEN_1498[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_19 <= _GEN_1499[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_20 <= _GEN_1500[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_21 <= _GEN_1501[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_22 <= _GEN_1502[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_23 <= _GEN_1503[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_24 <= _GEN_1504[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_25 <= _GEN_1505[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_26 <= _GEN_1506[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_27 <= _GEN_1507[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_28 <= _GEN_1508[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_29 <= _GEN_1509[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_30 <= _GEN_1510[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_31 <= _GEN_1511[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_32 <= _GEN_1512[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_33 <= _GEN_1513[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_34 <= _GEN_1514[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_35 <= _GEN_1515[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_36 <= _GEN_1516[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_37 <= _GEN_1517[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_38 <= _GEN_1518[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_39 <= _GEN_1519[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_40 <= _GEN_1520[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_41 <= _GEN_1521[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_42 <= _GEN_1522[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_43 <= _GEN_1523[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_44 <= _GEN_1524[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_45 <= _GEN_1525[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_46 <= _GEN_1526[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_47 <= _GEN_1527[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_48 <= _GEN_1528[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_49 <= _GEN_1529[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_50 <= _GEN_1530[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    a_aux_reg_r_51 <= _GEN_1531[105:0]; // @[BinaryDesigns2.scala 171:{30,30}]
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_0 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_0 <= 106'h1921fb54411744;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_1 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_1 <= b_aux_reg_r_0;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_2 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_2 <= b_aux_reg_r_1;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_3 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_3 <= b_aux_reg_r_2;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_4 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_4 <= b_aux_reg_r_3;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_5 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_5 <= b_aux_reg_r_4;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_6 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_6 <= b_aux_reg_r_5;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_7 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_7 <= b_aux_reg_r_6;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_8 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_8 <= b_aux_reg_r_7;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_9 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_9 <= b_aux_reg_r_8;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_10 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_10 <= b_aux_reg_r_9;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_11 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_11 <= b_aux_reg_r_10;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_12 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_12 <= b_aux_reg_r_11;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_13 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_13 <= b_aux_reg_r_12;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_14 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_14 <= b_aux_reg_r_13;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_15 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_15 <= b_aux_reg_r_14;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_16 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_16 <= b_aux_reg_r_15;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_17 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_17 <= b_aux_reg_r_16;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_18 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_18 <= b_aux_reg_r_17;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_19 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_19 <= b_aux_reg_r_18;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_20 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_20 <= b_aux_reg_r_19;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_21 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_21 <= b_aux_reg_r_20;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_22 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_22 <= b_aux_reg_r_21;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_23 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_23 <= b_aux_reg_r_22;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_24 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_24 <= b_aux_reg_r_23;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_25 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_25 <= b_aux_reg_r_24;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_26 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_26 <= b_aux_reg_r_25;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_27 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_27 <= b_aux_reg_r_26;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_28 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_28 <= b_aux_reg_r_27;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_29 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_29 <= b_aux_reg_r_28;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_30 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_30 <= b_aux_reg_r_29;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_31 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_31 <= b_aux_reg_r_30;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_32 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_32 <= b_aux_reg_r_31;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_33 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_33 <= b_aux_reg_r_32;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_34 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_34 <= b_aux_reg_r_33;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_35 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_35 <= b_aux_reg_r_34;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_36 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_36 <= b_aux_reg_r_35;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_37 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_37 <= b_aux_reg_r_36;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_38 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_38 <= b_aux_reg_r_37;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_39 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_39 <= b_aux_reg_r_38;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_40 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_40 <= b_aux_reg_r_39;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_41 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_41 <= b_aux_reg_r_40;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_42 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_42 <= b_aux_reg_r_41;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_43 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_43 <= b_aux_reg_r_42;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_44 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_44 <= b_aux_reg_r_43;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_45 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_45 <= b_aux_reg_r_44;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_46 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_46 <= b_aux_reg_r_45;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_47 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_47 <= b_aux_reg_r_46;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_48 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_48 <= b_aux_reg_r_47;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_49 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_49 <= b_aux_reg_r_48;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_50 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_50 <= b_aux_reg_r_49;
    end
    if (reset) begin // @[BinaryDesigns2.scala 176:30]
      b_aux_reg_r_51 <= 106'h0; // @[BinaryDesigns2.scala 176:30]
    end else begin
      b_aux_reg_r_51 <= b_aux_reg_r_50;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_1 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_1 <= _result_reg_r_1_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_2 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_2 <= _result_reg_r_2_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_3 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_3 <= _result_reg_r_3_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_4 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_4 <= _result_reg_r_4_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_5 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_5 <= _result_reg_r_5_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_6 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_6 <= _result_reg_r_6_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_7 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_7 <= _result_reg_r_7_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_8 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_8 <= _result_reg_r_8_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_9 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_9 <= _result_reg_r_9_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_10 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_10 <= _result_reg_r_10_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_11 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_11 <= _result_reg_r_11_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_12 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_12 <= _result_reg_r_12_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_13 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_13 <= _result_reg_r_13_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_14 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_14 <= _result_reg_r_14_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_15 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_15 <= _result_reg_r_15_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_16 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_16 <= _result_reg_r_16_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_17 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_17 <= _result_reg_r_17_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_18 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_18 <= _result_reg_r_18_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_19 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_19 <= _result_reg_r_19_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_20 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_20 <= _result_reg_r_20_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_21 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_21 <= _result_reg_r_21_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_22 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_22 <= _result_reg_r_22_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_23 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_23 <= _result_reg_r_23_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_24 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_24 <= _result_reg_r_24_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_25 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_25 <= _result_reg_r_25_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_26 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_26 <= _result_reg_r_26_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_27 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_27 <= _result_reg_r_27_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_28 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_28 <= _result_reg_r_28_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_29 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_29 <= _result_reg_r_29_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_30 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_30 <= _result_reg_r_30_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_31 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_31 <= _result_reg_r_31_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_32 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_32 <= _result_reg_r_32_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_33 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_33 <= _result_reg_r_33_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_34 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_34 <= _result_reg_r_34_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_35 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_35 <= _result_reg_r_35_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_36 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_36 <= _result_reg_r_36_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_37 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_37 <= _result_reg_r_37_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_38 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_38 <= _result_reg_r_38_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_39 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_39 <= _result_reg_r_39_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_40 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_40 <= _result_reg_r_40_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_41 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_41 <= _result_reg_r_41_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_42 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_42 <= _result_reg_r_42_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_43 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_43 <= _result_reg_r_43_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_44 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_44 <= _result_reg_r_44_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_45 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_45 <= _result_reg_r_45_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_46 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_46 <= _result_reg_r_46_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_47 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_47 <= _result_reg_r_47_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_48 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_48 <= _result_reg_r_48_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_49 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_49 <= _result_reg_r_49_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_50 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_50 <= _result_reg_r_50_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_51 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_51 <= _result_reg_r_51_T;
    end
    if (reset) begin // @[BinaryDesigns2.scala 181:31]
      result_reg_r_52 <= 106'h0; // @[BinaryDesigns2.scala 181:31]
    end else begin
      result_reg_r_52 <= _result_reg_r_52_T;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  a_aux_reg_r_0 = _RAND_0[105:0];
  _RAND_1 = {4{`RANDOM}};
  a_aux_reg_r_1 = _RAND_1[105:0];
  _RAND_2 = {4{`RANDOM}};
  a_aux_reg_r_2 = _RAND_2[105:0];
  _RAND_3 = {4{`RANDOM}};
  a_aux_reg_r_3 = _RAND_3[105:0];
  _RAND_4 = {4{`RANDOM}};
  a_aux_reg_r_4 = _RAND_4[105:0];
  _RAND_5 = {4{`RANDOM}};
  a_aux_reg_r_5 = _RAND_5[105:0];
  _RAND_6 = {4{`RANDOM}};
  a_aux_reg_r_6 = _RAND_6[105:0];
  _RAND_7 = {4{`RANDOM}};
  a_aux_reg_r_7 = _RAND_7[105:0];
  _RAND_8 = {4{`RANDOM}};
  a_aux_reg_r_8 = _RAND_8[105:0];
  _RAND_9 = {4{`RANDOM}};
  a_aux_reg_r_9 = _RAND_9[105:0];
  _RAND_10 = {4{`RANDOM}};
  a_aux_reg_r_10 = _RAND_10[105:0];
  _RAND_11 = {4{`RANDOM}};
  a_aux_reg_r_11 = _RAND_11[105:0];
  _RAND_12 = {4{`RANDOM}};
  a_aux_reg_r_12 = _RAND_12[105:0];
  _RAND_13 = {4{`RANDOM}};
  a_aux_reg_r_13 = _RAND_13[105:0];
  _RAND_14 = {4{`RANDOM}};
  a_aux_reg_r_14 = _RAND_14[105:0];
  _RAND_15 = {4{`RANDOM}};
  a_aux_reg_r_15 = _RAND_15[105:0];
  _RAND_16 = {4{`RANDOM}};
  a_aux_reg_r_16 = _RAND_16[105:0];
  _RAND_17 = {4{`RANDOM}};
  a_aux_reg_r_17 = _RAND_17[105:0];
  _RAND_18 = {4{`RANDOM}};
  a_aux_reg_r_18 = _RAND_18[105:0];
  _RAND_19 = {4{`RANDOM}};
  a_aux_reg_r_19 = _RAND_19[105:0];
  _RAND_20 = {4{`RANDOM}};
  a_aux_reg_r_20 = _RAND_20[105:0];
  _RAND_21 = {4{`RANDOM}};
  a_aux_reg_r_21 = _RAND_21[105:0];
  _RAND_22 = {4{`RANDOM}};
  a_aux_reg_r_22 = _RAND_22[105:0];
  _RAND_23 = {4{`RANDOM}};
  a_aux_reg_r_23 = _RAND_23[105:0];
  _RAND_24 = {4{`RANDOM}};
  a_aux_reg_r_24 = _RAND_24[105:0];
  _RAND_25 = {4{`RANDOM}};
  a_aux_reg_r_25 = _RAND_25[105:0];
  _RAND_26 = {4{`RANDOM}};
  a_aux_reg_r_26 = _RAND_26[105:0];
  _RAND_27 = {4{`RANDOM}};
  a_aux_reg_r_27 = _RAND_27[105:0];
  _RAND_28 = {4{`RANDOM}};
  a_aux_reg_r_28 = _RAND_28[105:0];
  _RAND_29 = {4{`RANDOM}};
  a_aux_reg_r_29 = _RAND_29[105:0];
  _RAND_30 = {4{`RANDOM}};
  a_aux_reg_r_30 = _RAND_30[105:0];
  _RAND_31 = {4{`RANDOM}};
  a_aux_reg_r_31 = _RAND_31[105:0];
  _RAND_32 = {4{`RANDOM}};
  a_aux_reg_r_32 = _RAND_32[105:0];
  _RAND_33 = {4{`RANDOM}};
  a_aux_reg_r_33 = _RAND_33[105:0];
  _RAND_34 = {4{`RANDOM}};
  a_aux_reg_r_34 = _RAND_34[105:0];
  _RAND_35 = {4{`RANDOM}};
  a_aux_reg_r_35 = _RAND_35[105:0];
  _RAND_36 = {4{`RANDOM}};
  a_aux_reg_r_36 = _RAND_36[105:0];
  _RAND_37 = {4{`RANDOM}};
  a_aux_reg_r_37 = _RAND_37[105:0];
  _RAND_38 = {4{`RANDOM}};
  a_aux_reg_r_38 = _RAND_38[105:0];
  _RAND_39 = {4{`RANDOM}};
  a_aux_reg_r_39 = _RAND_39[105:0];
  _RAND_40 = {4{`RANDOM}};
  a_aux_reg_r_40 = _RAND_40[105:0];
  _RAND_41 = {4{`RANDOM}};
  a_aux_reg_r_41 = _RAND_41[105:0];
  _RAND_42 = {4{`RANDOM}};
  a_aux_reg_r_42 = _RAND_42[105:0];
  _RAND_43 = {4{`RANDOM}};
  a_aux_reg_r_43 = _RAND_43[105:0];
  _RAND_44 = {4{`RANDOM}};
  a_aux_reg_r_44 = _RAND_44[105:0];
  _RAND_45 = {4{`RANDOM}};
  a_aux_reg_r_45 = _RAND_45[105:0];
  _RAND_46 = {4{`RANDOM}};
  a_aux_reg_r_46 = _RAND_46[105:0];
  _RAND_47 = {4{`RANDOM}};
  a_aux_reg_r_47 = _RAND_47[105:0];
  _RAND_48 = {4{`RANDOM}};
  a_aux_reg_r_48 = _RAND_48[105:0];
  _RAND_49 = {4{`RANDOM}};
  a_aux_reg_r_49 = _RAND_49[105:0];
  _RAND_50 = {4{`RANDOM}};
  a_aux_reg_r_50 = _RAND_50[105:0];
  _RAND_51 = {4{`RANDOM}};
  a_aux_reg_r_51 = _RAND_51[105:0];
  _RAND_52 = {4{`RANDOM}};
  b_aux_reg_r_0 = _RAND_52[105:0];
  _RAND_53 = {4{`RANDOM}};
  b_aux_reg_r_1 = _RAND_53[105:0];
  _RAND_54 = {4{`RANDOM}};
  b_aux_reg_r_2 = _RAND_54[105:0];
  _RAND_55 = {4{`RANDOM}};
  b_aux_reg_r_3 = _RAND_55[105:0];
  _RAND_56 = {4{`RANDOM}};
  b_aux_reg_r_4 = _RAND_56[105:0];
  _RAND_57 = {4{`RANDOM}};
  b_aux_reg_r_5 = _RAND_57[105:0];
  _RAND_58 = {4{`RANDOM}};
  b_aux_reg_r_6 = _RAND_58[105:0];
  _RAND_59 = {4{`RANDOM}};
  b_aux_reg_r_7 = _RAND_59[105:0];
  _RAND_60 = {4{`RANDOM}};
  b_aux_reg_r_8 = _RAND_60[105:0];
  _RAND_61 = {4{`RANDOM}};
  b_aux_reg_r_9 = _RAND_61[105:0];
  _RAND_62 = {4{`RANDOM}};
  b_aux_reg_r_10 = _RAND_62[105:0];
  _RAND_63 = {4{`RANDOM}};
  b_aux_reg_r_11 = _RAND_63[105:0];
  _RAND_64 = {4{`RANDOM}};
  b_aux_reg_r_12 = _RAND_64[105:0];
  _RAND_65 = {4{`RANDOM}};
  b_aux_reg_r_13 = _RAND_65[105:0];
  _RAND_66 = {4{`RANDOM}};
  b_aux_reg_r_14 = _RAND_66[105:0];
  _RAND_67 = {4{`RANDOM}};
  b_aux_reg_r_15 = _RAND_67[105:0];
  _RAND_68 = {4{`RANDOM}};
  b_aux_reg_r_16 = _RAND_68[105:0];
  _RAND_69 = {4{`RANDOM}};
  b_aux_reg_r_17 = _RAND_69[105:0];
  _RAND_70 = {4{`RANDOM}};
  b_aux_reg_r_18 = _RAND_70[105:0];
  _RAND_71 = {4{`RANDOM}};
  b_aux_reg_r_19 = _RAND_71[105:0];
  _RAND_72 = {4{`RANDOM}};
  b_aux_reg_r_20 = _RAND_72[105:0];
  _RAND_73 = {4{`RANDOM}};
  b_aux_reg_r_21 = _RAND_73[105:0];
  _RAND_74 = {4{`RANDOM}};
  b_aux_reg_r_22 = _RAND_74[105:0];
  _RAND_75 = {4{`RANDOM}};
  b_aux_reg_r_23 = _RAND_75[105:0];
  _RAND_76 = {4{`RANDOM}};
  b_aux_reg_r_24 = _RAND_76[105:0];
  _RAND_77 = {4{`RANDOM}};
  b_aux_reg_r_25 = _RAND_77[105:0];
  _RAND_78 = {4{`RANDOM}};
  b_aux_reg_r_26 = _RAND_78[105:0];
  _RAND_79 = {4{`RANDOM}};
  b_aux_reg_r_27 = _RAND_79[105:0];
  _RAND_80 = {4{`RANDOM}};
  b_aux_reg_r_28 = _RAND_80[105:0];
  _RAND_81 = {4{`RANDOM}};
  b_aux_reg_r_29 = _RAND_81[105:0];
  _RAND_82 = {4{`RANDOM}};
  b_aux_reg_r_30 = _RAND_82[105:0];
  _RAND_83 = {4{`RANDOM}};
  b_aux_reg_r_31 = _RAND_83[105:0];
  _RAND_84 = {4{`RANDOM}};
  b_aux_reg_r_32 = _RAND_84[105:0];
  _RAND_85 = {4{`RANDOM}};
  b_aux_reg_r_33 = _RAND_85[105:0];
  _RAND_86 = {4{`RANDOM}};
  b_aux_reg_r_34 = _RAND_86[105:0];
  _RAND_87 = {4{`RANDOM}};
  b_aux_reg_r_35 = _RAND_87[105:0];
  _RAND_88 = {4{`RANDOM}};
  b_aux_reg_r_36 = _RAND_88[105:0];
  _RAND_89 = {4{`RANDOM}};
  b_aux_reg_r_37 = _RAND_89[105:0];
  _RAND_90 = {4{`RANDOM}};
  b_aux_reg_r_38 = _RAND_90[105:0];
  _RAND_91 = {4{`RANDOM}};
  b_aux_reg_r_39 = _RAND_91[105:0];
  _RAND_92 = {4{`RANDOM}};
  b_aux_reg_r_40 = _RAND_92[105:0];
  _RAND_93 = {4{`RANDOM}};
  b_aux_reg_r_41 = _RAND_93[105:0];
  _RAND_94 = {4{`RANDOM}};
  b_aux_reg_r_42 = _RAND_94[105:0];
  _RAND_95 = {4{`RANDOM}};
  b_aux_reg_r_43 = _RAND_95[105:0];
  _RAND_96 = {4{`RANDOM}};
  b_aux_reg_r_44 = _RAND_96[105:0];
  _RAND_97 = {4{`RANDOM}};
  b_aux_reg_r_45 = _RAND_97[105:0];
  _RAND_98 = {4{`RANDOM}};
  b_aux_reg_r_46 = _RAND_98[105:0];
  _RAND_99 = {4{`RANDOM}};
  b_aux_reg_r_47 = _RAND_99[105:0];
  _RAND_100 = {4{`RANDOM}};
  b_aux_reg_r_48 = _RAND_100[105:0];
  _RAND_101 = {4{`RANDOM}};
  b_aux_reg_r_49 = _RAND_101[105:0];
  _RAND_102 = {4{`RANDOM}};
  b_aux_reg_r_50 = _RAND_102[105:0];
  _RAND_103 = {4{`RANDOM}};
  b_aux_reg_r_51 = _RAND_103[105:0];
  _RAND_104 = {4{`RANDOM}};
  result_reg_r_1 = _RAND_104[105:0];
  _RAND_105 = {4{`RANDOM}};
  result_reg_r_2 = _RAND_105[105:0];
  _RAND_106 = {4{`RANDOM}};
  result_reg_r_3 = _RAND_106[105:0];
  _RAND_107 = {4{`RANDOM}};
  result_reg_r_4 = _RAND_107[105:0];
  _RAND_108 = {4{`RANDOM}};
  result_reg_r_5 = _RAND_108[105:0];
  _RAND_109 = {4{`RANDOM}};
  result_reg_r_6 = _RAND_109[105:0];
  _RAND_110 = {4{`RANDOM}};
  result_reg_r_7 = _RAND_110[105:0];
  _RAND_111 = {4{`RANDOM}};
  result_reg_r_8 = _RAND_111[105:0];
  _RAND_112 = {4{`RANDOM}};
  result_reg_r_9 = _RAND_112[105:0];
  _RAND_113 = {4{`RANDOM}};
  result_reg_r_10 = _RAND_113[105:0];
  _RAND_114 = {4{`RANDOM}};
  result_reg_r_11 = _RAND_114[105:0];
  _RAND_115 = {4{`RANDOM}};
  result_reg_r_12 = _RAND_115[105:0];
  _RAND_116 = {4{`RANDOM}};
  result_reg_r_13 = _RAND_116[105:0];
  _RAND_117 = {4{`RANDOM}};
  result_reg_r_14 = _RAND_117[105:0];
  _RAND_118 = {4{`RANDOM}};
  result_reg_r_15 = _RAND_118[105:0];
  _RAND_119 = {4{`RANDOM}};
  result_reg_r_16 = _RAND_119[105:0];
  _RAND_120 = {4{`RANDOM}};
  result_reg_r_17 = _RAND_120[105:0];
  _RAND_121 = {4{`RANDOM}};
  result_reg_r_18 = _RAND_121[105:0];
  _RAND_122 = {4{`RANDOM}};
  result_reg_r_19 = _RAND_122[105:0];
  _RAND_123 = {4{`RANDOM}};
  result_reg_r_20 = _RAND_123[105:0];
  _RAND_124 = {4{`RANDOM}};
  result_reg_r_21 = _RAND_124[105:0];
  _RAND_125 = {4{`RANDOM}};
  result_reg_r_22 = _RAND_125[105:0];
  _RAND_126 = {4{`RANDOM}};
  result_reg_r_23 = _RAND_126[105:0];
  _RAND_127 = {4{`RANDOM}};
  result_reg_r_24 = _RAND_127[105:0];
  _RAND_128 = {4{`RANDOM}};
  result_reg_r_25 = _RAND_128[105:0];
  _RAND_129 = {4{`RANDOM}};
  result_reg_r_26 = _RAND_129[105:0];
  _RAND_130 = {4{`RANDOM}};
  result_reg_r_27 = _RAND_130[105:0];
  _RAND_131 = {4{`RANDOM}};
  result_reg_r_28 = _RAND_131[105:0];
  _RAND_132 = {4{`RANDOM}};
  result_reg_r_29 = _RAND_132[105:0];
  _RAND_133 = {4{`RANDOM}};
  result_reg_r_30 = _RAND_133[105:0];
  _RAND_134 = {4{`RANDOM}};
  result_reg_r_31 = _RAND_134[105:0];
  _RAND_135 = {4{`RANDOM}};
  result_reg_r_32 = _RAND_135[105:0];
  _RAND_136 = {4{`RANDOM}};
  result_reg_r_33 = _RAND_136[105:0];
  _RAND_137 = {4{`RANDOM}};
  result_reg_r_34 = _RAND_137[105:0];
  _RAND_138 = {4{`RANDOM}};
  result_reg_r_35 = _RAND_138[105:0];
  _RAND_139 = {4{`RANDOM}};
  result_reg_r_36 = _RAND_139[105:0];
  _RAND_140 = {4{`RANDOM}};
  result_reg_r_37 = _RAND_140[105:0];
  _RAND_141 = {4{`RANDOM}};
  result_reg_r_38 = _RAND_141[105:0];
  _RAND_142 = {4{`RANDOM}};
  result_reg_r_39 = _RAND_142[105:0];
  _RAND_143 = {4{`RANDOM}};
  result_reg_r_40 = _RAND_143[105:0];
  _RAND_144 = {4{`RANDOM}};
  result_reg_r_41 = _RAND_144[105:0];
  _RAND_145 = {4{`RANDOM}};
  result_reg_r_42 = _RAND_145[105:0];
  _RAND_146 = {4{`RANDOM}};
  result_reg_r_43 = _RAND_146[105:0];
  _RAND_147 = {4{`RANDOM}};
  result_reg_r_44 = _RAND_147[105:0];
  _RAND_148 = {4{`RANDOM}};
  result_reg_r_45 = _RAND_148[105:0];
  _RAND_149 = {4{`RANDOM}};
  result_reg_r_46 = _RAND_149[105:0];
  _RAND_150 = {4{`RANDOM}};
  result_reg_r_47 = _RAND_150[105:0];
  _RAND_151 = {4{`RANDOM}};
  result_reg_r_48 = _RAND_151[105:0];
  _RAND_152 = {4{`RANDOM}};
  result_reg_r_49 = _RAND_152[105:0];
  _RAND_153 = {4{`RANDOM}};
  result_reg_r_50 = _RAND_153[105:0];
  _RAND_154 = {4{`RANDOM}};
  result_reg_r_51 = _RAND_154[105:0];
  _RAND_155 = {4{`RANDOM}};
  result_reg_r_52 = _RAND_155[105:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
