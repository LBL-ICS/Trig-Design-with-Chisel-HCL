module CLZ128(
  input  [127:0] io_in,
  output [6:0]   io_out
);
  wire [127:0] _ax_T = io_in & 128'hffffffffffffffff0000000000000000; // @[FixedPoint.scala 211:20]
  wire  _ax_T_1 = _ax_T == 128'h0; // @[FixedPoint.scala 211:29]
  wire [191:0] _ax_T_2 = {io_in, 64'h0}; // @[FixedPoint.scala 211:41]
  wire [191:0] ax = _ax_T == 128'h0 ? _ax_T_2 : {{64'd0}, io_in}; // @[FixedPoint.scala 211:15]
  wire [191:0] _bx_T = ax & 192'hffffffff000000000000000000000000; // @[FixedPoint.scala 212:20]
  wire  _bx_T_1 = _bx_T == 192'h0; // @[FixedPoint.scala 212:29]
  wire [223:0] _bx_T_2 = {ax, 32'h0}; // @[FixedPoint.scala 212:41]
  wire [223:0] bx = _bx_T == 192'h0 ? _bx_T_2 : {{32'd0}, ax}; // @[FixedPoint.scala 212:15]
  wire [223:0] _cx_T = bx & 224'hffff0000000000000000000000000000; // @[FixedPoint.scala 213:20]
  wire  _cx_T_1 = _cx_T == 224'h0; // @[FixedPoint.scala 213:29]
  wire [239:0] _cx_T_2 = {bx, 16'h0}; // @[FixedPoint.scala 213:41]
  wire [239:0] cx = _cx_T == 224'h0 ? _cx_T_2 : {{16'd0}, bx}; // @[FixedPoint.scala 213:15]
  wire [239:0] _dx_T = cx & 240'hff000000000000000000000000000000; // @[FixedPoint.scala 214:20]
  wire  _dx_T_1 = _dx_T == 240'h0; // @[FixedPoint.scala 214:29]
  wire [247:0] _dx_T_2 = {cx, 8'h0}; // @[FixedPoint.scala 214:41]
  wire [247:0] dx = _dx_T == 240'h0 ? _dx_T_2 : {{8'd0}, cx}; // @[FixedPoint.scala 214:15]
  wire [247:0] _ex_T = dx & 248'hf0000000000000000000000000000000; // @[FixedPoint.scala 215:20]
  wire  _ex_T_1 = _ex_T == 248'h0; // @[FixedPoint.scala 215:29]
  wire [251:0] _ex_T_2 = {dx, 4'h0}; // @[FixedPoint.scala 215:41]
  wire [251:0] ex = _ex_T == 248'h0 ? _ex_T_2 : {{4'd0}, dx}; // @[FixedPoint.scala 215:15]
  wire [251:0] _fx_T = ex & 252'hc0000000000000000000000000000000; // @[FixedPoint.scala 216:20]
  wire  _fx_T_1 = _fx_T == 252'h0; // @[FixedPoint.scala 216:29]
  wire [253:0] _fx_T_2 = {ex, 2'h0}; // @[FixedPoint.scala 216:41]
  wire [253:0] fx = _fx_T == 252'h0 ? _fx_T_2 : {{2'd0}, ex}; // @[FixedPoint.scala 216:15]
  wire [5:0] _io_out_T_16 = {_ax_T_1,_bx_T_1,_cx_T_1,_dx_T_1,_ex_T_1,_fx_T_1}; // @[FixedPoint.scala 223:28]
  wire [253:0] _io_out_T_17 = fx & 254'h80000000000000000000000000000000; // @[FixedPoint.scala 225:10]
  wire  _io_out_T_18 = _io_out_T_17 == 254'h0; // @[FixedPoint.scala 225:19]
  assign io_out = {_io_out_T_16,_io_out_T_18}; // @[FixedPoint.scala 224:29]
endmodule
