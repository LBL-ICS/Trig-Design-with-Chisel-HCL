module FP_divider_bw128(
  input          clock,
  input          reset,
  input  [127:0] io_in_a,
  output [127:0] io_out_s
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
`endif // RANDOMIZE_REG_INIT
  wire [14:0] postProcess_exp_subtractor_io_in_a; // @[FloatingPointDesigns2.scala 499:44]
  wire [14:0] postProcess_exp_subtractor_io_in_b; // @[FloatingPointDesigns2.scala 499:44]
  wire [14:0] postProcess_exp_subtractor_io_out_s; // @[FloatingPointDesigns2.scala 499:44]
  wire  postProcess_exp_subtractor_io_out_c; // @[FloatingPointDesigns2.scala 499:44]
  wire  divider_BW226_v3_clock; // @[FloatingPointDesigns2.scala 504:30]
  wire  divider_BW226_v3_reset; // @[FloatingPointDesigns2.scala 504:30]
  wire [225:0] divider_BW226_v3_io_in_a; // @[FloatingPointDesigns2.scala 504:30]
  wire [225:0] divider_BW226_v3_io_out_s; // @[FloatingPointDesigns2.scala 504:30]
  wire [14:0] _GEN_0 = io_in_a[126:112] < 15'h1 ? 15'h1 : io_in_a[126:112]; // @[FloatingPointDesigns2.scala 472:49 473:19 475:19]
  wire [111:0] frac_wire_0 = io_in_a[111:0]; // @[FloatingPointDesigns2.scala 487:28]
  wire [112:0] whole_frac_wire_0 = {1'h1,frac_wire_0}; // @[FloatingPointDesigns2.scala 492:31]
  reg  carry_flag_r; // @[Reg.scala 16:16]
  reg  carry_flag_r_1; // @[Reg.scala 16:16]
  reg  carry_flag_r_2; // @[Reg.scala 16:16]
  reg  carry_flag_r_3; // @[Reg.scala 16:16]
  reg  carry_flag_r_4; // @[Reg.scala 16:16]
  reg  carry_flag_r_5; // @[Reg.scala 16:16]
  reg  carry_flag_r_6; // @[Reg.scala 16:16]
  reg  carry_flag_r_7; // @[Reg.scala 16:16]
  reg  carry_flag_r_8; // @[Reg.scala 16:16]
  reg  carry_flag_r_9; // @[Reg.scala 16:16]
  reg  carry_flag_r_10; // @[Reg.scala 16:16]
  reg  carry_flag_r_11; // @[Reg.scala 16:16]
  reg  carry_flag_r_12; // @[Reg.scala 16:16]
  reg  carry_flag_r_13; // @[Reg.scala 16:16]
  reg  carry_flag_r_14; // @[Reg.scala 16:16]
  reg  carry_flag_r_15; // @[Reg.scala 16:16]
  reg  carry_flag_r_16; // @[Reg.scala 16:16]
  reg  carry_flag_r_17; // @[Reg.scala 16:16]
  reg  carry_flag_r_18; // @[Reg.scala 16:16]
  reg  carry_flag_r_19; // @[Reg.scala 16:16]
  reg  carry_flag_r_20; // @[Reg.scala 16:16]
  reg  carry_flag_r_21; // @[Reg.scala 16:16]
  reg  carry_flag_r_22; // @[Reg.scala 16:16]
  reg  carry_flag_r_23; // @[Reg.scala 16:16]
  reg  carry_flag_r_24; // @[Reg.scala 16:16]
  reg  carry_flag_r_25; // @[Reg.scala 16:16]
  reg  carry_flag_r_26; // @[Reg.scala 16:16]
  reg  carry_flag_r_27; // @[Reg.scala 16:16]
  reg  carry_flag_r_28; // @[Reg.scala 16:16]
  reg  carry_flag_r_29; // @[Reg.scala 16:16]
  reg  carry_flag_r_30; // @[Reg.scala 16:16]
  reg  carry_flag_r_31; // @[Reg.scala 16:16]
  reg  carry_flag_r_32; // @[Reg.scala 16:16]
  reg  carry_flag_r_33; // @[Reg.scala 16:16]
  reg  carry_flag_r_34; // @[Reg.scala 16:16]
  reg  carry_flag_r_35; // @[Reg.scala 16:16]
  reg  carry_flag_r_36; // @[Reg.scala 16:16]
  reg  carry_flag_r_37; // @[Reg.scala 16:16]
  reg  carry_flag_r_38; // @[Reg.scala 16:16]
  reg  carry_flag_r_39; // @[Reg.scala 16:16]
  reg  carry_flag_r_40; // @[Reg.scala 16:16]
  reg  carry_flag_r_41; // @[Reg.scala 16:16]
  reg  carry_flag_r_42; // @[Reg.scala 16:16]
  reg  carry_flag_r_43; // @[Reg.scala 16:16]
  reg  carry_flag_r_44; // @[Reg.scala 16:16]
  reg  carry_flag_r_45; // @[Reg.scala 16:16]
  reg  carry_flag_r_46; // @[Reg.scala 16:16]
  reg  carry_flag_r_47; // @[Reg.scala 16:16]
  reg  carry_flag_r_48; // @[Reg.scala 16:16]
  reg  carry_flag_r_49; // @[Reg.scala 16:16]
  reg  carry_flag_r_50; // @[Reg.scala 16:16]
  reg  carry_flag_r_51; // @[Reg.scala 16:16]
  reg  carry_flag_r_52; // @[Reg.scala 16:16]
  reg  carry_flag_r_53; // @[Reg.scala 16:16]
  reg  carry_flag_r_54; // @[Reg.scala 16:16]
  reg  carry_flag_r_55; // @[Reg.scala 16:16]
  reg  carry_flag_r_56; // @[Reg.scala 16:16]
  reg  carry_flag_r_57; // @[Reg.scala 16:16]
  reg  carry_flag_r_58; // @[Reg.scala 16:16]
  reg  carry_flag_r_59; // @[Reg.scala 16:16]
  reg  carry_flag_r_60; // @[Reg.scala 16:16]
  reg  carry_flag_r_61; // @[Reg.scala 16:16]
  reg  carry_flag_r_62; // @[Reg.scala 16:16]
  reg  carry_flag_r_63; // @[Reg.scala 16:16]
  reg  carry_flag_r_64; // @[Reg.scala 16:16]
  reg  carry_flag_r_65; // @[Reg.scala 16:16]
  reg  carry_flag_r_66; // @[Reg.scala 16:16]
  reg  carry_flag_r_67; // @[Reg.scala 16:16]
  reg  carry_flag_r_68; // @[Reg.scala 16:16]
  reg  carry_flag_r_69; // @[Reg.scala 16:16]
  reg  carry_flag_r_70; // @[Reg.scala 16:16]
  reg  carry_flag_r_71; // @[Reg.scala 16:16]
  reg  carry_flag_r_72; // @[Reg.scala 16:16]
  reg  carry_flag_r_73; // @[Reg.scala 16:16]
  reg  carry_flag_r_74; // @[Reg.scala 16:16]
  reg  carry_flag_r_75; // @[Reg.scala 16:16]
  reg  carry_flag_r_76; // @[Reg.scala 16:16]
  reg  carry_flag_r_77; // @[Reg.scala 16:16]
  reg  carry_flag_r_78; // @[Reg.scala 16:16]
  reg  carry_flag_r_79; // @[Reg.scala 16:16]
  reg  carry_flag_r_80; // @[Reg.scala 16:16]
  reg  carry_flag_r_81; // @[Reg.scala 16:16]
  reg  carry_flag_r_82; // @[Reg.scala 16:16]
  reg  carry_flag_r_83; // @[Reg.scala 16:16]
  reg  carry_flag_r_84; // @[Reg.scala 16:16]
  reg  carry_flag_r_85; // @[Reg.scala 16:16]
  reg  carry_flag_r_86; // @[Reg.scala 16:16]
  reg  carry_flag_r_87; // @[Reg.scala 16:16]
  reg  carry_flag_r_88; // @[Reg.scala 16:16]
  reg  carry_flag_r_89; // @[Reg.scala 16:16]
  reg  carry_flag_r_90; // @[Reg.scala 16:16]
  reg  carry_flag_r_91; // @[Reg.scala 16:16]
  reg  carry_flag_r_92; // @[Reg.scala 16:16]
  reg  carry_flag_r_93; // @[Reg.scala 16:16]
  reg  carry_flag_r_94; // @[Reg.scala 16:16]
  reg  carry_flag_r_95; // @[Reg.scala 16:16]
  reg  carry_flag_r_96; // @[Reg.scala 16:16]
  reg  carry_flag_r_97; // @[Reg.scala 16:16]
  reg  carry_flag_r_98; // @[Reg.scala 16:16]
  reg  carry_flag_r_99; // @[Reg.scala 16:16]
  reg  carry_flag_r_100; // @[Reg.scala 16:16]
  reg  carry_flag_r_101; // @[Reg.scala 16:16]
  reg  carry_flag_r_102; // @[Reg.scala 16:16]
  reg  carry_flag_r_103; // @[Reg.scala 16:16]
  reg  carry_flag_r_104; // @[Reg.scala 16:16]
  reg  carry_flag_r_105; // @[Reg.scala 16:16]
  reg  carry_flag_r_106; // @[Reg.scala 16:16]
  reg  carry_flag_r_107; // @[Reg.scala 16:16]
  reg  carry_flag_r_108; // @[Reg.scala 16:16]
  reg  carry_flag_r_109; // @[Reg.scala 16:16]
  reg  carry_flag_r_110; // @[Reg.scala 16:16]
  reg  carry_flag_r_111; // @[Reg.scala 16:16]
  reg  carry_flag; // @[Reg.scala 16:16]
  wire  msb_check = divider_BW226_v3_io_out_s[113]; // @[FloatingPointDesigns2.scala 513:39]
  reg [14:0] exp_sum_r; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_1; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_2; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_3; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_4; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_5; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_6; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_7; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_8; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_9; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_10; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_11; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_12; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_13; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_14; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_15; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_16; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_17; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_18; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_19; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_20; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_21; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_22; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_23; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_24; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_25; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_26; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_27; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_28; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_29; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_30; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_31; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_32; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_33; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_34; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_35; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_36; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_37; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_38; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_39; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_40; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_41; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_42; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_43; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_44; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_45; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_46; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_47; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_48; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_49; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_50; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_51; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_52; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_53; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_54; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_55; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_56; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_57; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_58; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_59; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_60; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_61; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_62; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_63; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_64; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_65; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_66; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_67; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_68; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_69; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_70; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_71; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_72; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_73; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_74; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_75; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_76; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_77; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_78; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_79; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_80; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_81; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_82; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_83; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_84; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_85; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_86; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_87; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_88; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_89; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_90; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_91; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_92; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_93; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_94; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_95; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_96; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_97; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_98; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_99; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_100; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_101; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_102; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_103; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_104; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_105; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_106; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_107; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_108; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_109; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_110; // @[Reg.scala 16:16]
  reg [14:0] exp_sum_r_111; // @[Reg.scala 16:16]
  reg [14:0] exp_sum; // @[Reg.scala 16:16]
  reg  new_sign_reg_r; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_1; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_2; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_3; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_4; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_5; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_6; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_7; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_8; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_9; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_10; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_11; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_12; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_13; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_14; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_15; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_16; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_17; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_18; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_19; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_20; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_21; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_22; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_23; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_24; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_25; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_26; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_27; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_28; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_29; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_30; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_31; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_32; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_33; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_34; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_35; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_36; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_37; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_38; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_39; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_40; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_41; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_42; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_43; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_44; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_45; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_46; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_47; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_48; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_49; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_50; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_51; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_52; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_53; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_54; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_55; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_56; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_57; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_58; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_59; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_60; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_61; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_62; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_63; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_64; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_65; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_66; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_67; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_68; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_69; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_70; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_71; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_72; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_73; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_74; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_75; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_76; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_77; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_78; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_79; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_80; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_81; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_82; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_83; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_84; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_85; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_86; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_87; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_88; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_89; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_90; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_91; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_92; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_93; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_94; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_95; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_96; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_97; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_98; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_99; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_100; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_101; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_102; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_103; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_104; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_105; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_106; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_107; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_108; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_109; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_110; // @[Reg.scala 16:16]
  reg  new_sign_reg_r_111; // @[Reg.scala 16:16]
  reg  new_sign_reg; // @[Reg.scala 16:16]
  wire  _u_flag_reg_T_1 = ~msb_check; // @[FloatingPointDesigns2.scala 519:64]
  wire [14:0] _GEN_456 = {{14'd0}, _u_flag_reg_T_1}; // @[FloatingPointDesigns2.scala 519:60]
  wire [15:0] _u_flag_reg_T_2 = exp_sum - _GEN_456; // @[FloatingPointDesigns2.scala 519:60]
  wire  o_flag_reg = carry_flag | _u_flag_reg_T_2 < 16'h1; // @[FloatingPointDesigns2.scala 520:47]
  wire [14:0] _out_exp_T_1 = exp_sum - 15'h1; // @[FloatingPointDesigns2.scala 526:109]
  wire [14:0] _out_exp_T_2 = msb_check ? exp_sum : _out_exp_T_1; // @[FloatingPointDesigns2.scala 526:72]
  wire [14:0] out_exp = o_flag_reg ? 15'h1 : _out_exp_T_2; // @[FloatingPointDesigns2.scala 526:47]
  wire [111:0] _out_frac_T_2 = msb_check ? divider_BW226_v3_io_out_s[112:1] : divider_BW226_v3_io_out_s[111:0]; // @[FloatingPointDesigns2.scala 527:74]
  wire [111:0] out_frac = o_flag_reg ? 112'h0 : _out_frac_T_2; // @[FloatingPointDesigns2.scala 527:49]
  wire [15:0] _io_out_s_T = {new_sign_reg,out_exp}; // @[FloatingPointDesigns2.scala 528:26]
  full_subtractor postProcess_exp_subtractor ( // @[FloatingPointDesigns2.scala 499:44]
    .io_in_a(postProcess_exp_subtractor_io_in_a),
    .io_in_b(postProcess_exp_subtractor_io_in_b),
    .io_out_s(postProcess_exp_subtractor_io_out_s),
    .io_out_c(postProcess_exp_subtractor_io_out_c)
  );
  divider_BW226_v3 divider_BW226_v3 ( // @[FloatingPointDesigns2.scala 504:30]
    .clock(divider_BW226_v3_clock),
    .reset(divider_BW226_v3_reset),
    .io_in_a(divider_BW226_v3_io_in_a),
    .io_out_s(divider_BW226_v3_io_out_s)
  );
  assign io_out_s = {_io_out_s_T,out_frac}; // @[FloatingPointDesigns2.scala 528:37]
  assign postProcess_exp_subtractor_io_in_a = io_in_a[126:112] > 15'h7ffe ? 15'h7ffe : _GEN_0; // @[FloatingPointDesigns2.scala 470:47 471:19]
  assign postProcess_exp_subtractor_io_in_b = 15'h4001 - 15'h3fff; // @[FloatingPointDesigns2.scala 501:55]
  assign divider_BW226_v3_clock = clock;
  assign divider_BW226_v3_reset = reset;
  assign divider_BW226_v3_io_in_a = {whole_frac_wire_0,113'h0}; // @[FloatingPointDesigns2.scala 508:45]
  always @(posedge clock) begin
    carry_flag_r <= postProcess_exp_subtractor_io_out_c; // @[FloatingPointDesigns2.scala 512:72]
    carry_flag_r_1 <= carry_flag_r; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_2 <= carry_flag_r_1; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_3 <= carry_flag_r_2; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_4 <= carry_flag_r_3; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_5 <= carry_flag_r_4; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_6 <= carry_flag_r_5; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_7 <= carry_flag_r_6; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_8 <= carry_flag_r_7; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_9 <= carry_flag_r_8; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_10 <= carry_flag_r_9; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_11 <= carry_flag_r_10; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_12 <= carry_flag_r_11; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_13 <= carry_flag_r_12; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_14 <= carry_flag_r_13; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_15 <= carry_flag_r_14; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_16 <= carry_flag_r_15; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_17 <= carry_flag_r_16; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_18 <= carry_flag_r_17; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_19 <= carry_flag_r_18; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_20 <= carry_flag_r_19; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_21 <= carry_flag_r_20; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_22 <= carry_flag_r_21; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_23 <= carry_flag_r_22; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_24 <= carry_flag_r_23; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_25 <= carry_flag_r_24; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_26 <= carry_flag_r_25; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_27 <= carry_flag_r_26; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_28 <= carry_flag_r_27; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_29 <= carry_flag_r_28; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_30 <= carry_flag_r_29; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_31 <= carry_flag_r_30; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_32 <= carry_flag_r_31; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_33 <= carry_flag_r_32; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_34 <= carry_flag_r_33; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_35 <= carry_flag_r_34; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_36 <= carry_flag_r_35; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_37 <= carry_flag_r_36; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_38 <= carry_flag_r_37; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_39 <= carry_flag_r_38; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_40 <= carry_flag_r_39; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_41 <= carry_flag_r_40; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_42 <= carry_flag_r_41; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_43 <= carry_flag_r_42; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_44 <= carry_flag_r_43; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_45 <= carry_flag_r_44; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_46 <= carry_flag_r_45; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_47 <= carry_flag_r_46; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_48 <= carry_flag_r_47; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_49 <= carry_flag_r_48; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_50 <= carry_flag_r_49; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_51 <= carry_flag_r_50; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_52 <= carry_flag_r_51; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_53 <= carry_flag_r_52; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_54 <= carry_flag_r_53; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_55 <= carry_flag_r_54; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_56 <= carry_flag_r_55; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_57 <= carry_flag_r_56; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_58 <= carry_flag_r_57; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_59 <= carry_flag_r_58; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_60 <= carry_flag_r_59; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_61 <= carry_flag_r_60; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_62 <= carry_flag_r_61; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_63 <= carry_flag_r_62; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_64 <= carry_flag_r_63; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_65 <= carry_flag_r_64; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_66 <= carry_flag_r_65; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_67 <= carry_flag_r_66; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_68 <= carry_flag_r_67; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_69 <= carry_flag_r_68; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_70 <= carry_flag_r_69; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_71 <= carry_flag_r_70; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_72 <= carry_flag_r_71; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_73 <= carry_flag_r_72; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_74 <= carry_flag_r_73; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_75 <= carry_flag_r_74; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_76 <= carry_flag_r_75; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_77 <= carry_flag_r_76; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_78 <= carry_flag_r_77; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_79 <= carry_flag_r_78; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_80 <= carry_flag_r_79; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_81 <= carry_flag_r_80; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_82 <= carry_flag_r_81; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_83 <= carry_flag_r_82; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_84 <= carry_flag_r_83; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_85 <= carry_flag_r_84; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_86 <= carry_flag_r_85; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_87 <= carry_flag_r_86; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_88 <= carry_flag_r_87; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_89 <= carry_flag_r_88; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_90 <= carry_flag_r_89; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_91 <= carry_flag_r_90; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_92 <= carry_flag_r_91; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_93 <= carry_flag_r_92; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_94 <= carry_flag_r_93; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_95 <= carry_flag_r_94; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_96 <= carry_flag_r_95; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_97 <= carry_flag_r_96; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_98 <= carry_flag_r_97; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_99 <= carry_flag_r_98; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_100 <= carry_flag_r_99; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_101 <= carry_flag_r_100; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_102 <= carry_flag_r_101; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_103 <= carry_flag_r_102; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_104 <= carry_flag_r_103; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_105 <= carry_flag_r_104; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_106 <= carry_flag_r_105; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_107 <= carry_flag_r_106; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_108 <= carry_flag_r_107; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_109 <= carry_flag_r_108; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_110 <= carry_flag_r_109; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag_r_111 <= carry_flag_r_110; // @[Reg.scala 16:16 17:{18,22}]
    carry_flag <= carry_flag_r_111; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r <= postProcess_exp_subtractor_io_out_s; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_1 <= exp_sum_r; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_2 <= exp_sum_r_1; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_3 <= exp_sum_r_2; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_4 <= exp_sum_r_3; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_5 <= exp_sum_r_4; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_6 <= exp_sum_r_5; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_7 <= exp_sum_r_6; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_8 <= exp_sum_r_7; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_9 <= exp_sum_r_8; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_10 <= exp_sum_r_9; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_11 <= exp_sum_r_10; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_12 <= exp_sum_r_11; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_13 <= exp_sum_r_12; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_14 <= exp_sum_r_13; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_15 <= exp_sum_r_14; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_16 <= exp_sum_r_15; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_17 <= exp_sum_r_16; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_18 <= exp_sum_r_17; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_19 <= exp_sum_r_18; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_20 <= exp_sum_r_19; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_21 <= exp_sum_r_20; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_22 <= exp_sum_r_21; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_23 <= exp_sum_r_22; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_24 <= exp_sum_r_23; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_25 <= exp_sum_r_24; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_26 <= exp_sum_r_25; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_27 <= exp_sum_r_26; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_28 <= exp_sum_r_27; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_29 <= exp_sum_r_28; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_30 <= exp_sum_r_29; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_31 <= exp_sum_r_30; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_32 <= exp_sum_r_31; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_33 <= exp_sum_r_32; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_34 <= exp_sum_r_33; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_35 <= exp_sum_r_34; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_36 <= exp_sum_r_35; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_37 <= exp_sum_r_36; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_38 <= exp_sum_r_37; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_39 <= exp_sum_r_38; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_40 <= exp_sum_r_39; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_41 <= exp_sum_r_40; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_42 <= exp_sum_r_41; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_43 <= exp_sum_r_42; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_44 <= exp_sum_r_43; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_45 <= exp_sum_r_44; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_46 <= exp_sum_r_45; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_47 <= exp_sum_r_46; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_48 <= exp_sum_r_47; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_49 <= exp_sum_r_48; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_50 <= exp_sum_r_49; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_51 <= exp_sum_r_50; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_52 <= exp_sum_r_51; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_53 <= exp_sum_r_52; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_54 <= exp_sum_r_53; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_55 <= exp_sum_r_54; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_56 <= exp_sum_r_55; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_57 <= exp_sum_r_56; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_58 <= exp_sum_r_57; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_59 <= exp_sum_r_58; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_60 <= exp_sum_r_59; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_61 <= exp_sum_r_60; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_62 <= exp_sum_r_61; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_63 <= exp_sum_r_62; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_64 <= exp_sum_r_63; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_65 <= exp_sum_r_64; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_66 <= exp_sum_r_65; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_67 <= exp_sum_r_66; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_68 <= exp_sum_r_67; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_69 <= exp_sum_r_68; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_70 <= exp_sum_r_69; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_71 <= exp_sum_r_70; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_72 <= exp_sum_r_71; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_73 <= exp_sum_r_72; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_74 <= exp_sum_r_73; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_75 <= exp_sum_r_74; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_76 <= exp_sum_r_75; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_77 <= exp_sum_r_76; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_78 <= exp_sum_r_77; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_79 <= exp_sum_r_78; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_80 <= exp_sum_r_79; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_81 <= exp_sum_r_80; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_82 <= exp_sum_r_81; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_83 <= exp_sum_r_82; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_84 <= exp_sum_r_83; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_85 <= exp_sum_r_84; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_86 <= exp_sum_r_85; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_87 <= exp_sum_r_86; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_88 <= exp_sum_r_87; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_89 <= exp_sum_r_88; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_90 <= exp_sum_r_89; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_91 <= exp_sum_r_90; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_92 <= exp_sum_r_91; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_93 <= exp_sum_r_92; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_94 <= exp_sum_r_93; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_95 <= exp_sum_r_94; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_96 <= exp_sum_r_95; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_97 <= exp_sum_r_96; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_98 <= exp_sum_r_97; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_99 <= exp_sum_r_98; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_100 <= exp_sum_r_99; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_101 <= exp_sum_r_100; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_102 <= exp_sum_r_101; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_103 <= exp_sum_r_102; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_104 <= exp_sum_r_103; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_105 <= exp_sum_r_104; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_106 <= exp_sum_r_105; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_107 <= exp_sum_r_106; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_108 <= exp_sum_r_107; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_109 <= exp_sum_r_108; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_110 <= exp_sum_r_109; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum_r_111 <= exp_sum_r_110; // @[Reg.scala 16:16 17:{18,22}]
    exp_sum <= exp_sum_r_111; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r <= io_in_a[127]; // @[FloatingPointDesigns2.scala 465:28]
    new_sign_reg_r_1 <= new_sign_reg_r; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_2 <= new_sign_reg_r_1; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_3 <= new_sign_reg_r_2; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_4 <= new_sign_reg_r_3; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_5 <= new_sign_reg_r_4; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_6 <= new_sign_reg_r_5; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_7 <= new_sign_reg_r_6; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_8 <= new_sign_reg_r_7; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_9 <= new_sign_reg_r_8; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_10 <= new_sign_reg_r_9; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_11 <= new_sign_reg_r_10; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_12 <= new_sign_reg_r_11; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_13 <= new_sign_reg_r_12; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_14 <= new_sign_reg_r_13; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_15 <= new_sign_reg_r_14; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_16 <= new_sign_reg_r_15; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_17 <= new_sign_reg_r_16; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_18 <= new_sign_reg_r_17; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_19 <= new_sign_reg_r_18; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_20 <= new_sign_reg_r_19; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_21 <= new_sign_reg_r_20; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_22 <= new_sign_reg_r_21; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_23 <= new_sign_reg_r_22; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_24 <= new_sign_reg_r_23; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_25 <= new_sign_reg_r_24; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_26 <= new_sign_reg_r_25; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_27 <= new_sign_reg_r_26; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_28 <= new_sign_reg_r_27; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_29 <= new_sign_reg_r_28; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_30 <= new_sign_reg_r_29; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_31 <= new_sign_reg_r_30; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_32 <= new_sign_reg_r_31; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_33 <= new_sign_reg_r_32; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_34 <= new_sign_reg_r_33; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_35 <= new_sign_reg_r_34; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_36 <= new_sign_reg_r_35; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_37 <= new_sign_reg_r_36; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_38 <= new_sign_reg_r_37; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_39 <= new_sign_reg_r_38; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_40 <= new_sign_reg_r_39; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_41 <= new_sign_reg_r_40; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_42 <= new_sign_reg_r_41; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_43 <= new_sign_reg_r_42; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_44 <= new_sign_reg_r_43; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_45 <= new_sign_reg_r_44; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_46 <= new_sign_reg_r_45; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_47 <= new_sign_reg_r_46; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_48 <= new_sign_reg_r_47; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_49 <= new_sign_reg_r_48; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_50 <= new_sign_reg_r_49; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_51 <= new_sign_reg_r_50; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_52 <= new_sign_reg_r_51; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_53 <= new_sign_reg_r_52; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_54 <= new_sign_reg_r_53; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_55 <= new_sign_reg_r_54; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_56 <= new_sign_reg_r_55; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_57 <= new_sign_reg_r_56; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_58 <= new_sign_reg_r_57; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_59 <= new_sign_reg_r_58; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_60 <= new_sign_reg_r_59; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_61 <= new_sign_reg_r_60; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_62 <= new_sign_reg_r_61; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_63 <= new_sign_reg_r_62; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_64 <= new_sign_reg_r_63; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_65 <= new_sign_reg_r_64; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_66 <= new_sign_reg_r_65; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_67 <= new_sign_reg_r_66; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_68 <= new_sign_reg_r_67; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_69 <= new_sign_reg_r_68; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_70 <= new_sign_reg_r_69; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_71 <= new_sign_reg_r_70; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_72 <= new_sign_reg_r_71; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_73 <= new_sign_reg_r_72; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_74 <= new_sign_reg_r_73; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_75 <= new_sign_reg_r_74; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_76 <= new_sign_reg_r_75; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_77 <= new_sign_reg_r_76; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_78 <= new_sign_reg_r_77; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_79 <= new_sign_reg_r_78; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_80 <= new_sign_reg_r_79; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_81 <= new_sign_reg_r_80; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_82 <= new_sign_reg_r_81; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_83 <= new_sign_reg_r_82; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_84 <= new_sign_reg_r_83; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_85 <= new_sign_reg_r_84; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_86 <= new_sign_reg_r_85; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_87 <= new_sign_reg_r_86; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_88 <= new_sign_reg_r_87; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_89 <= new_sign_reg_r_88; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_90 <= new_sign_reg_r_89; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_91 <= new_sign_reg_r_90; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_92 <= new_sign_reg_r_91; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_93 <= new_sign_reg_r_92; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_94 <= new_sign_reg_r_93; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_95 <= new_sign_reg_r_94; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_96 <= new_sign_reg_r_95; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_97 <= new_sign_reg_r_96; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_98 <= new_sign_reg_r_97; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_99 <= new_sign_reg_r_98; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_100 <= new_sign_reg_r_99; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_101 <= new_sign_reg_r_100; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_102 <= new_sign_reg_r_101; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_103 <= new_sign_reg_r_102; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_104 <= new_sign_reg_r_103; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_105 <= new_sign_reg_r_104; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_106 <= new_sign_reg_r_105; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_107 <= new_sign_reg_r_106; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_108 <= new_sign_reg_r_107; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_109 <= new_sign_reg_r_108; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_110 <= new_sign_reg_r_109; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg_r_111 <= new_sign_reg_r_110; // @[Reg.scala 16:16 17:{18,22}]
    new_sign_reg <= new_sign_reg_r_111; // @[Reg.scala 16:16 17:{18,22}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  carry_flag_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  carry_flag_r_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  carry_flag_r_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  carry_flag_r_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  carry_flag_r_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  carry_flag_r_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  carry_flag_r_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  carry_flag_r_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  carry_flag_r_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  carry_flag_r_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  carry_flag_r_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  carry_flag_r_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  carry_flag_r_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  carry_flag_r_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  carry_flag_r_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  carry_flag_r_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  carry_flag_r_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  carry_flag_r_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  carry_flag_r_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  carry_flag_r_19 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  carry_flag_r_20 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  carry_flag_r_21 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  carry_flag_r_22 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  carry_flag_r_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  carry_flag_r_24 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  carry_flag_r_25 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  carry_flag_r_26 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  carry_flag_r_27 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  carry_flag_r_28 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  carry_flag_r_29 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  carry_flag_r_30 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  carry_flag_r_31 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  carry_flag_r_32 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  carry_flag_r_33 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  carry_flag_r_34 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  carry_flag_r_35 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  carry_flag_r_36 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  carry_flag_r_37 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  carry_flag_r_38 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  carry_flag_r_39 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  carry_flag_r_40 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  carry_flag_r_41 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  carry_flag_r_42 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  carry_flag_r_43 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  carry_flag_r_44 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  carry_flag_r_45 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  carry_flag_r_46 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  carry_flag_r_47 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  carry_flag_r_48 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  carry_flag_r_49 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  carry_flag_r_50 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  carry_flag_r_51 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  carry_flag_r_52 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  carry_flag_r_53 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  carry_flag_r_54 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  carry_flag_r_55 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  carry_flag_r_56 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  carry_flag_r_57 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  carry_flag_r_58 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  carry_flag_r_59 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  carry_flag_r_60 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  carry_flag_r_61 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  carry_flag_r_62 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  carry_flag_r_63 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  carry_flag_r_64 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  carry_flag_r_65 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  carry_flag_r_66 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  carry_flag_r_67 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  carry_flag_r_68 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  carry_flag_r_69 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  carry_flag_r_70 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  carry_flag_r_71 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  carry_flag_r_72 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  carry_flag_r_73 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  carry_flag_r_74 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  carry_flag_r_75 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  carry_flag_r_76 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  carry_flag_r_77 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  carry_flag_r_78 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  carry_flag_r_79 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  carry_flag_r_80 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  carry_flag_r_81 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  carry_flag_r_82 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  carry_flag_r_83 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  carry_flag_r_84 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  carry_flag_r_85 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  carry_flag_r_86 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  carry_flag_r_87 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  carry_flag_r_88 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  carry_flag_r_89 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  carry_flag_r_90 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  carry_flag_r_91 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  carry_flag_r_92 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  carry_flag_r_93 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  carry_flag_r_94 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  carry_flag_r_95 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  carry_flag_r_96 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  carry_flag_r_97 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  carry_flag_r_98 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  carry_flag_r_99 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  carry_flag_r_100 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  carry_flag_r_101 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  carry_flag_r_102 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  carry_flag_r_103 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  carry_flag_r_104 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  carry_flag_r_105 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  carry_flag_r_106 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  carry_flag_r_107 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  carry_flag_r_108 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  carry_flag_r_109 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  carry_flag_r_110 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  carry_flag_r_111 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  carry_flag = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  exp_sum_r = _RAND_113[14:0];
  _RAND_114 = {1{`RANDOM}};
  exp_sum_r_1 = _RAND_114[14:0];
  _RAND_115 = {1{`RANDOM}};
  exp_sum_r_2 = _RAND_115[14:0];
  _RAND_116 = {1{`RANDOM}};
  exp_sum_r_3 = _RAND_116[14:0];
  _RAND_117 = {1{`RANDOM}};
  exp_sum_r_4 = _RAND_117[14:0];
  _RAND_118 = {1{`RANDOM}};
  exp_sum_r_5 = _RAND_118[14:0];
  _RAND_119 = {1{`RANDOM}};
  exp_sum_r_6 = _RAND_119[14:0];
  _RAND_120 = {1{`RANDOM}};
  exp_sum_r_7 = _RAND_120[14:0];
  _RAND_121 = {1{`RANDOM}};
  exp_sum_r_8 = _RAND_121[14:0];
  _RAND_122 = {1{`RANDOM}};
  exp_sum_r_9 = _RAND_122[14:0];
  _RAND_123 = {1{`RANDOM}};
  exp_sum_r_10 = _RAND_123[14:0];
  _RAND_124 = {1{`RANDOM}};
  exp_sum_r_11 = _RAND_124[14:0];
  _RAND_125 = {1{`RANDOM}};
  exp_sum_r_12 = _RAND_125[14:0];
  _RAND_126 = {1{`RANDOM}};
  exp_sum_r_13 = _RAND_126[14:0];
  _RAND_127 = {1{`RANDOM}};
  exp_sum_r_14 = _RAND_127[14:0];
  _RAND_128 = {1{`RANDOM}};
  exp_sum_r_15 = _RAND_128[14:0];
  _RAND_129 = {1{`RANDOM}};
  exp_sum_r_16 = _RAND_129[14:0];
  _RAND_130 = {1{`RANDOM}};
  exp_sum_r_17 = _RAND_130[14:0];
  _RAND_131 = {1{`RANDOM}};
  exp_sum_r_18 = _RAND_131[14:0];
  _RAND_132 = {1{`RANDOM}};
  exp_sum_r_19 = _RAND_132[14:0];
  _RAND_133 = {1{`RANDOM}};
  exp_sum_r_20 = _RAND_133[14:0];
  _RAND_134 = {1{`RANDOM}};
  exp_sum_r_21 = _RAND_134[14:0];
  _RAND_135 = {1{`RANDOM}};
  exp_sum_r_22 = _RAND_135[14:0];
  _RAND_136 = {1{`RANDOM}};
  exp_sum_r_23 = _RAND_136[14:0];
  _RAND_137 = {1{`RANDOM}};
  exp_sum_r_24 = _RAND_137[14:0];
  _RAND_138 = {1{`RANDOM}};
  exp_sum_r_25 = _RAND_138[14:0];
  _RAND_139 = {1{`RANDOM}};
  exp_sum_r_26 = _RAND_139[14:0];
  _RAND_140 = {1{`RANDOM}};
  exp_sum_r_27 = _RAND_140[14:0];
  _RAND_141 = {1{`RANDOM}};
  exp_sum_r_28 = _RAND_141[14:0];
  _RAND_142 = {1{`RANDOM}};
  exp_sum_r_29 = _RAND_142[14:0];
  _RAND_143 = {1{`RANDOM}};
  exp_sum_r_30 = _RAND_143[14:0];
  _RAND_144 = {1{`RANDOM}};
  exp_sum_r_31 = _RAND_144[14:0];
  _RAND_145 = {1{`RANDOM}};
  exp_sum_r_32 = _RAND_145[14:0];
  _RAND_146 = {1{`RANDOM}};
  exp_sum_r_33 = _RAND_146[14:0];
  _RAND_147 = {1{`RANDOM}};
  exp_sum_r_34 = _RAND_147[14:0];
  _RAND_148 = {1{`RANDOM}};
  exp_sum_r_35 = _RAND_148[14:0];
  _RAND_149 = {1{`RANDOM}};
  exp_sum_r_36 = _RAND_149[14:0];
  _RAND_150 = {1{`RANDOM}};
  exp_sum_r_37 = _RAND_150[14:0];
  _RAND_151 = {1{`RANDOM}};
  exp_sum_r_38 = _RAND_151[14:0];
  _RAND_152 = {1{`RANDOM}};
  exp_sum_r_39 = _RAND_152[14:0];
  _RAND_153 = {1{`RANDOM}};
  exp_sum_r_40 = _RAND_153[14:0];
  _RAND_154 = {1{`RANDOM}};
  exp_sum_r_41 = _RAND_154[14:0];
  _RAND_155 = {1{`RANDOM}};
  exp_sum_r_42 = _RAND_155[14:0];
  _RAND_156 = {1{`RANDOM}};
  exp_sum_r_43 = _RAND_156[14:0];
  _RAND_157 = {1{`RANDOM}};
  exp_sum_r_44 = _RAND_157[14:0];
  _RAND_158 = {1{`RANDOM}};
  exp_sum_r_45 = _RAND_158[14:0];
  _RAND_159 = {1{`RANDOM}};
  exp_sum_r_46 = _RAND_159[14:0];
  _RAND_160 = {1{`RANDOM}};
  exp_sum_r_47 = _RAND_160[14:0];
  _RAND_161 = {1{`RANDOM}};
  exp_sum_r_48 = _RAND_161[14:0];
  _RAND_162 = {1{`RANDOM}};
  exp_sum_r_49 = _RAND_162[14:0];
  _RAND_163 = {1{`RANDOM}};
  exp_sum_r_50 = _RAND_163[14:0];
  _RAND_164 = {1{`RANDOM}};
  exp_sum_r_51 = _RAND_164[14:0];
  _RAND_165 = {1{`RANDOM}};
  exp_sum_r_52 = _RAND_165[14:0];
  _RAND_166 = {1{`RANDOM}};
  exp_sum_r_53 = _RAND_166[14:0];
  _RAND_167 = {1{`RANDOM}};
  exp_sum_r_54 = _RAND_167[14:0];
  _RAND_168 = {1{`RANDOM}};
  exp_sum_r_55 = _RAND_168[14:0];
  _RAND_169 = {1{`RANDOM}};
  exp_sum_r_56 = _RAND_169[14:0];
  _RAND_170 = {1{`RANDOM}};
  exp_sum_r_57 = _RAND_170[14:0];
  _RAND_171 = {1{`RANDOM}};
  exp_sum_r_58 = _RAND_171[14:0];
  _RAND_172 = {1{`RANDOM}};
  exp_sum_r_59 = _RAND_172[14:0];
  _RAND_173 = {1{`RANDOM}};
  exp_sum_r_60 = _RAND_173[14:0];
  _RAND_174 = {1{`RANDOM}};
  exp_sum_r_61 = _RAND_174[14:0];
  _RAND_175 = {1{`RANDOM}};
  exp_sum_r_62 = _RAND_175[14:0];
  _RAND_176 = {1{`RANDOM}};
  exp_sum_r_63 = _RAND_176[14:0];
  _RAND_177 = {1{`RANDOM}};
  exp_sum_r_64 = _RAND_177[14:0];
  _RAND_178 = {1{`RANDOM}};
  exp_sum_r_65 = _RAND_178[14:0];
  _RAND_179 = {1{`RANDOM}};
  exp_sum_r_66 = _RAND_179[14:0];
  _RAND_180 = {1{`RANDOM}};
  exp_sum_r_67 = _RAND_180[14:0];
  _RAND_181 = {1{`RANDOM}};
  exp_sum_r_68 = _RAND_181[14:0];
  _RAND_182 = {1{`RANDOM}};
  exp_sum_r_69 = _RAND_182[14:0];
  _RAND_183 = {1{`RANDOM}};
  exp_sum_r_70 = _RAND_183[14:0];
  _RAND_184 = {1{`RANDOM}};
  exp_sum_r_71 = _RAND_184[14:0];
  _RAND_185 = {1{`RANDOM}};
  exp_sum_r_72 = _RAND_185[14:0];
  _RAND_186 = {1{`RANDOM}};
  exp_sum_r_73 = _RAND_186[14:0];
  _RAND_187 = {1{`RANDOM}};
  exp_sum_r_74 = _RAND_187[14:0];
  _RAND_188 = {1{`RANDOM}};
  exp_sum_r_75 = _RAND_188[14:0];
  _RAND_189 = {1{`RANDOM}};
  exp_sum_r_76 = _RAND_189[14:0];
  _RAND_190 = {1{`RANDOM}};
  exp_sum_r_77 = _RAND_190[14:0];
  _RAND_191 = {1{`RANDOM}};
  exp_sum_r_78 = _RAND_191[14:0];
  _RAND_192 = {1{`RANDOM}};
  exp_sum_r_79 = _RAND_192[14:0];
  _RAND_193 = {1{`RANDOM}};
  exp_sum_r_80 = _RAND_193[14:0];
  _RAND_194 = {1{`RANDOM}};
  exp_sum_r_81 = _RAND_194[14:0];
  _RAND_195 = {1{`RANDOM}};
  exp_sum_r_82 = _RAND_195[14:0];
  _RAND_196 = {1{`RANDOM}};
  exp_sum_r_83 = _RAND_196[14:0];
  _RAND_197 = {1{`RANDOM}};
  exp_sum_r_84 = _RAND_197[14:0];
  _RAND_198 = {1{`RANDOM}};
  exp_sum_r_85 = _RAND_198[14:0];
  _RAND_199 = {1{`RANDOM}};
  exp_sum_r_86 = _RAND_199[14:0];
  _RAND_200 = {1{`RANDOM}};
  exp_sum_r_87 = _RAND_200[14:0];
  _RAND_201 = {1{`RANDOM}};
  exp_sum_r_88 = _RAND_201[14:0];
  _RAND_202 = {1{`RANDOM}};
  exp_sum_r_89 = _RAND_202[14:0];
  _RAND_203 = {1{`RANDOM}};
  exp_sum_r_90 = _RAND_203[14:0];
  _RAND_204 = {1{`RANDOM}};
  exp_sum_r_91 = _RAND_204[14:0];
  _RAND_205 = {1{`RANDOM}};
  exp_sum_r_92 = _RAND_205[14:0];
  _RAND_206 = {1{`RANDOM}};
  exp_sum_r_93 = _RAND_206[14:0];
  _RAND_207 = {1{`RANDOM}};
  exp_sum_r_94 = _RAND_207[14:0];
  _RAND_208 = {1{`RANDOM}};
  exp_sum_r_95 = _RAND_208[14:0];
  _RAND_209 = {1{`RANDOM}};
  exp_sum_r_96 = _RAND_209[14:0];
  _RAND_210 = {1{`RANDOM}};
  exp_sum_r_97 = _RAND_210[14:0];
  _RAND_211 = {1{`RANDOM}};
  exp_sum_r_98 = _RAND_211[14:0];
  _RAND_212 = {1{`RANDOM}};
  exp_sum_r_99 = _RAND_212[14:0];
  _RAND_213 = {1{`RANDOM}};
  exp_sum_r_100 = _RAND_213[14:0];
  _RAND_214 = {1{`RANDOM}};
  exp_sum_r_101 = _RAND_214[14:0];
  _RAND_215 = {1{`RANDOM}};
  exp_sum_r_102 = _RAND_215[14:0];
  _RAND_216 = {1{`RANDOM}};
  exp_sum_r_103 = _RAND_216[14:0];
  _RAND_217 = {1{`RANDOM}};
  exp_sum_r_104 = _RAND_217[14:0];
  _RAND_218 = {1{`RANDOM}};
  exp_sum_r_105 = _RAND_218[14:0];
  _RAND_219 = {1{`RANDOM}};
  exp_sum_r_106 = _RAND_219[14:0];
  _RAND_220 = {1{`RANDOM}};
  exp_sum_r_107 = _RAND_220[14:0];
  _RAND_221 = {1{`RANDOM}};
  exp_sum_r_108 = _RAND_221[14:0];
  _RAND_222 = {1{`RANDOM}};
  exp_sum_r_109 = _RAND_222[14:0];
  _RAND_223 = {1{`RANDOM}};
  exp_sum_r_110 = _RAND_223[14:0];
  _RAND_224 = {1{`RANDOM}};
  exp_sum_r_111 = _RAND_224[14:0];
  _RAND_225 = {1{`RANDOM}};
  exp_sum = _RAND_225[14:0];
  _RAND_226 = {1{`RANDOM}};
  new_sign_reg_r = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  new_sign_reg_r_1 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  new_sign_reg_r_2 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  new_sign_reg_r_3 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  new_sign_reg_r_4 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  new_sign_reg_r_5 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  new_sign_reg_r_6 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  new_sign_reg_r_7 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  new_sign_reg_r_8 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  new_sign_reg_r_9 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  new_sign_reg_r_10 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  new_sign_reg_r_11 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  new_sign_reg_r_12 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  new_sign_reg_r_13 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  new_sign_reg_r_14 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  new_sign_reg_r_15 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  new_sign_reg_r_16 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  new_sign_reg_r_17 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  new_sign_reg_r_18 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  new_sign_reg_r_19 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  new_sign_reg_r_20 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  new_sign_reg_r_21 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  new_sign_reg_r_22 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  new_sign_reg_r_23 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  new_sign_reg_r_24 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  new_sign_reg_r_25 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  new_sign_reg_r_26 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  new_sign_reg_r_27 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  new_sign_reg_r_28 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  new_sign_reg_r_29 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  new_sign_reg_r_30 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  new_sign_reg_r_31 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  new_sign_reg_r_32 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  new_sign_reg_r_33 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  new_sign_reg_r_34 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  new_sign_reg_r_35 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  new_sign_reg_r_36 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  new_sign_reg_r_37 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  new_sign_reg_r_38 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  new_sign_reg_r_39 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  new_sign_reg_r_40 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  new_sign_reg_r_41 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  new_sign_reg_r_42 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  new_sign_reg_r_43 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  new_sign_reg_r_44 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  new_sign_reg_r_45 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  new_sign_reg_r_46 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  new_sign_reg_r_47 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  new_sign_reg_r_48 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  new_sign_reg_r_49 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  new_sign_reg_r_50 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  new_sign_reg_r_51 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  new_sign_reg_r_52 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  new_sign_reg_r_53 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  new_sign_reg_r_54 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  new_sign_reg_r_55 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  new_sign_reg_r_56 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  new_sign_reg_r_57 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  new_sign_reg_r_58 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  new_sign_reg_r_59 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  new_sign_reg_r_60 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  new_sign_reg_r_61 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  new_sign_reg_r_62 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  new_sign_reg_r_63 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  new_sign_reg_r_64 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  new_sign_reg_r_65 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  new_sign_reg_r_66 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  new_sign_reg_r_67 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  new_sign_reg_r_68 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  new_sign_reg_r_69 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  new_sign_reg_r_70 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  new_sign_reg_r_71 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  new_sign_reg_r_72 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  new_sign_reg_r_73 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  new_sign_reg_r_74 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  new_sign_reg_r_75 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  new_sign_reg_r_76 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  new_sign_reg_r_77 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  new_sign_reg_r_78 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  new_sign_reg_r_79 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  new_sign_reg_r_80 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  new_sign_reg_r_81 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  new_sign_reg_r_82 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  new_sign_reg_r_83 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  new_sign_reg_r_84 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  new_sign_reg_r_85 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  new_sign_reg_r_86 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  new_sign_reg_r_87 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  new_sign_reg_r_88 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  new_sign_reg_r_89 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  new_sign_reg_r_90 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  new_sign_reg_r_91 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  new_sign_reg_r_92 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  new_sign_reg_r_93 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  new_sign_reg_r_94 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  new_sign_reg_r_95 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  new_sign_reg_r_96 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  new_sign_reg_r_97 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  new_sign_reg_r_98 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  new_sign_reg_r_99 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  new_sign_reg_r_100 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  new_sign_reg_r_101 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  new_sign_reg_r_102 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  new_sign_reg_r_103 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  new_sign_reg_r_104 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  new_sign_reg_r_105 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  new_sign_reg_r_106 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  new_sign_reg_r_107 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  new_sign_reg_r_108 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  new_sign_reg_r_109 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  new_sign_reg_r_110 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  new_sign_reg_r_111 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  new_sign_reg = _RAND_338[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
