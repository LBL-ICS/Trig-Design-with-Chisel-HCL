module leadingOneDetector(
  input  [111:0] io_in,
  output [6:0]   io_out
);
  wire [1:0] _hotValue_T = io_in[1] ? 2'h2 : 2'h1; // @[Mux.scala 47:70]
  wire [1:0] _hotValue_T_1 = io_in[2] ? 2'h3 : _hotValue_T; // @[Mux.scala 47:70]
  wire [2:0] _hotValue_T_2 = io_in[3] ? 3'h4 : {{1'd0}, _hotValue_T_1}; // @[Mux.scala 47:70]
  wire [2:0] _hotValue_T_3 = io_in[4] ? 3'h5 : _hotValue_T_2; // @[Mux.scala 47:70]
  wire [2:0] _hotValue_T_4 = io_in[5] ? 3'h6 : _hotValue_T_3; // @[Mux.scala 47:70]
  wire [2:0] _hotValue_T_5 = io_in[6] ? 3'h7 : _hotValue_T_4; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_6 = io_in[7] ? 4'h8 : {{1'd0}, _hotValue_T_5}; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_7 = io_in[8] ? 4'h9 : _hotValue_T_6; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_8 = io_in[9] ? 4'ha : _hotValue_T_7; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_9 = io_in[10] ? 4'hb : _hotValue_T_8; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_10 = io_in[11] ? 4'hc : _hotValue_T_9; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_11 = io_in[12] ? 4'hd : _hotValue_T_10; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_12 = io_in[13] ? 4'he : _hotValue_T_11; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_13 = io_in[14] ? 4'hf : _hotValue_T_12; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_14 = io_in[15] ? 5'h10 : {{1'd0}, _hotValue_T_13}; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_15 = io_in[16] ? 5'h11 : _hotValue_T_14; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_16 = io_in[17] ? 5'h12 : _hotValue_T_15; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_17 = io_in[18] ? 5'h13 : _hotValue_T_16; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_18 = io_in[19] ? 5'h14 : _hotValue_T_17; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_19 = io_in[20] ? 5'h15 : _hotValue_T_18; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_20 = io_in[21] ? 5'h16 : _hotValue_T_19; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_21 = io_in[22] ? 5'h17 : _hotValue_T_20; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_22 = io_in[23] ? 5'h18 : _hotValue_T_21; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_23 = io_in[24] ? 5'h19 : _hotValue_T_22; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_24 = io_in[25] ? 5'h1a : _hotValue_T_23; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_25 = io_in[26] ? 5'h1b : _hotValue_T_24; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_26 = io_in[27] ? 5'h1c : _hotValue_T_25; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_27 = io_in[28] ? 5'h1d : _hotValue_T_26; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_28 = io_in[29] ? 5'h1e : _hotValue_T_27; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_29 = io_in[30] ? 5'h1f : _hotValue_T_28; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_30 = io_in[31] ? 6'h20 : {{1'd0}, _hotValue_T_29}; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_31 = io_in[32] ? 6'h21 : _hotValue_T_30; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_32 = io_in[33] ? 6'h22 : _hotValue_T_31; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_33 = io_in[34] ? 6'h23 : _hotValue_T_32; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_34 = io_in[35] ? 6'h24 : _hotValue_T_33; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_35 = io_in[36] ? 6'h25 : _hotValue_T_34; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_36 = io_in[37] ? 6'h26 : _hotValue_T_35; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_37 = io_in[38] ? 6'h27 : _hotValue_T_36; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_38 = io_in[39] ? 6'h28 : _hotValue_T_37; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_39 = io_in[40] ? 6'h29 : _hotValue_T_38; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_40 = io_in[41] ? 6'h2a : _hotValue_T_39; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_41 = io_in[42] ? 6'h2b : _hotValue_T_40; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_42 = io_in[43] ? 6'h2c : _hotValue_T_41; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_43 = io_in[44] ? 6'h2d : _hotValue_T_42; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_44 = io_in[45] ? 6'h2e : _hotValue_T_43; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_45 = io_in[46] ? 6'h2f : _hotValue_T_44; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_46 = io_in[47] ? 6'h30 : _hotValue_T_45; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_47 = io_in[48] ? 6'h31 : _hotValue_T_46; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_48 = io_in[49] ? 6'h32 : _hotValue_T_47; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_49 = io_in[50] ? 6'h33 : _hotValue_T_48; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_50 = io_in[51] ? 6'h34 : _hotValue_T_49; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_51 = io_in[52] ? 6'h35 : _hotValue_T_50; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_52 = io_in[53] ? 6'h36 : _hotValue_T_51; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_53 = io_in[54] ? 6'h37 : _hotValue_T_52; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_54 = io_in[55] ? 6'h38 : _hotValue_T_53; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_55 = io_in[56] ? 6'h39 : _hotValue_T_54; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_56 = io_in[57] ? 6'h3a : _hotValue_T_55; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_57 = io_in[58] ? 6'h3b : _hotValue_T_56; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_58 = io_in[59] ? 6'h3c : _hotValue_T_57; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_59 = io_in[60] ? 6'h3d : _hotValue_T_58; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_60 = io_in[61] ? 6'h3e : _hotValue_T_59; // @[Mux.scala 47:70]
  wire [5:0] _hotValue_T_61 = io_in[62] ? 6'h3f : _hotValue_T_60; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_62 = io_in[63] ? 7'h40 : {{1'd0}, _hotValue_T_61}; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_63 = io_in[64] ? 7'h41 : _hotValue_T_62; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_64 = io_in[65] ? 7'h42 : _hotValue_T_63; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_65 = io_in[66] ? 7'h43 : _hotValue_T_64; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_66 = io_in[67] ? 7'h44 : _hotValue_T_65; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_67 = io_in[68] ? 7'h45 : _hotValue_T_66; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_68 = io_in[69] ? 7'h46 : _hotValue_T_67; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_69 = io_in[70] ? 7'h47 : _hotValue_T_68; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_70 = io_in[71] ? 7'h48 : _hotValue_T_69; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_71 = io_in[72] ? 7'h49 : _hotValue_T_70; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_72 = io_in[73] ? 7'h4a : _hotValue_T_71; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_73 = io_in[74] ? 7'h4b : _hotValue_T_72; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_74 = io_in[75] ? 7'h4c : _hotValue_T_73; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_75 = io_in[76] ? 7'h4d : _hotValue_T_74; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_76 = io_in[77] ? 7'h4e : _hotValue_T_75; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_77 = io_in[78] ? 7'h4f : _hotValue_T_76; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_78 = io_in[79] ? 7'h50 : _hotValue_T_77; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_79 = io_in[80] ? 7'h51 : _hotValue_T_78; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_80 = io_in[81] ? 7'h52 : _hotValue_T_79; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_81 = io_in[82] ? 7'h53 : _hotValue_T_80; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_82 = io_in[83] ? 7'h54 : _hotValue_T_81; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_83 = io_in[84] ? 7'h55 : _hotValue_T_82; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_84 = io_in[85] ? 7'h56 : _hotValue_T_83; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_85 = io_in[86] ? 7'h57 : _hotValue_T_84; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_86 = io_in[87] ? 7'h58 : _hotValue_T_85; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_87 = io_in[88] ? 7'h59 : _hotValue_T_86; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_88 = io_in[89] ? 7'h5a : _hotValue_T_87; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_89 = io_in[90] ? 7'h5b : _hotValue_T_88; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_90 = io_in[91] ? 7'h5c : _hotValue_T_89; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_91 = io_in[92] ? 7'h5d : _hotValue_T_90; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_92 = io_in[93] ? 7'h5e : _hotValue_T_91; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_93 = io_in[94] ? 7'h5f : _hotValue_T_92; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_94 = io_in[95] ? 7'h60 : _hotValue_T_93; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_95 = io_in[96] ? 7'h61 : _hotValue_T_94; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_96 = io_in[97] ? 7'h62 : _hotValue_T_95; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_97 = io_in[98] ? 7'h63 : _hotValue_T_96; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_98 = io_in[99] ? 7'h64 : _hotValue_T_97; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_99 = io_in[100] ? 7'h65 : _hotValue_T_98; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_100 = io_in[101] ? 7'h66 : _hotValue_T_99; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_101 = io_in[102] ? 7'h67 : _hotValue_T_100; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_102 = io_in[103] ? 7'h68 : _hotValue_T_101; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_103 = io_in[104] ? 7'h69 : _hotValue_T_102; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_104 = io_in[105] ? 7'h6a : _hotValue_T_103; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_105 = io_in[106] ? 7'h6b : _hotValue_T_104; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_106 = io_in[107] ? 7'h6c : _hotValue_T_105; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_107 = io_in[108] ? 7'h6d : _hotValue_T_106; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_108 = io_in[109] ? 7'h6e : _hotValue_T_107; // @[Mux.scala 47:70]
  wire [6:0] _hotValue_T_109 = io_in[110] ? 7'h6f : _hotValue_T_108; // @[Mux.scala 47:70]
  assign io_out = io_in[111] ? 7'h70 : _hotValue_T_109; // @[Mux.scala 47:70]
endmodule
